library verilog;
use verilog.vl_types.all;
entity proj1_testbench is
end proj1_testbench;
