
module mips_core ( clk, rst, cop_dout, din, ins_i, iack_o, cop_addr_o, 
        cop_data_o, cop_mem_ctl_o, addr_o, dout, pc_o, wr_en_o );
  input [31:0] cop_dout;
  input [31:0] din;
  input [31:0] ins_i;
  output [31:0] cop_addr_o;
  output [31:0] cop_data_o;
  output [3:0] cop_mem_ctl_o;
  output [31:0] addr_o;
  output [31:0] dout;
  output [31:0] pc_o;
  output [3:0] wr_en_o;
  input clk, rst;
  output iack_o;
  wire   NET1375, NET767, NET457, \MEM_CTL/BUS629[1] , \MEM_CTL/BUS629[0] ,
         \iRF_stage/BUS3236[4] , \iRF_stage/BUS3236[3] ,
         \iRF_stage/BUS3236[2] , \iRF_stage/BUS3236[1] ,
         \iRF_stage/BUS3236[0] , \iRF_stage/BUS3237[4] ,
         \iRF_stage/BUS3237[3] , \iRF_stage/BUS3237[2] ,
         \iRF_stage/BUS3237[1] , \iRF_stage/BUS3237[0] ,
         \iexec_stage/BUS2332[31] , \iexec_stage/BUS2332[30] ,
         \iexec_stage/BUS2332[29] , \iexec_stage/BUS2332[28] ,
         \iexec_stage/BUS2332[27] , \iexec_stage/BUS2332[26] ,
         \iexec_stage/BUS2332[25] , \iexec_stage/BUS2332[24] ,
         \iexec_stage/BUS2332[23] , \iexec_stage/BUS2332[22] ,
         \iexec_stage/BUS2332[21] , \iexec_stage/BUS2332[20] ,
         \iexec_stage/BUS2332[19] , \iexec_stage/BUS2332[18] ,
         \iexec_stage/BUS2332[17] , \iexec_stage/BUS2332[16] ,
         \iexec_stage/BUS2332[15] , \iexec_stage/BUS2332[14] ,
         \iexec_stage/BUS2332[13] , \iexec_stage/BUS2332[12] ,
         \iexec_stage/BUS2332[11] , \iexec_stage/BUS2332[10] ,
         \iexec_stage/BUS2332[9] , \iexec_stage/BUS2332[8] ,
         \iexec_stage/BUS2332[7] , \iexec_stage/BUS2332[6] ,
         \iexec_stage/BUS2332[5] , \iexec_stage/BUS2332[4] ,
         \iexec_stage/BUS2332[3] , \iexec_stage/BUS2332[2] ,
         \iexec_stage/BUS2332[1] , \iexec_stage/BUS2332[0] ,
         \iexec_stage/BUS2446[31] , \iexec_stage/BUS2446[30] ,
         \iexec_stage/BUS2446[29] , \iexec_stage/BUS2446[28] ,
         \iexec_stage/BUS2446[27] , \iexec_stage/BUS2446[26] ,
         \iexec_stage/BUS2446[25] , \iexec_stage/BUS2446[24] ,
         \iexec_stage/BUS2446[23] , \iexec_stage/BUS2446[22] ,
         \iexec_stage/BUS2446[21] , \iexec_stage/BUS2446[20] ,
         \iexec_stage/BUS2446[19] , \iexec_stage/BUS2446[18] ,
         \iexec_stage/BUS2446[17] , \iexec_stage/BUS2446[16] ,
         \iexec_stage/BUS2446[15] , \iexec_stage/BUS2446[14] ,
         \iexec_stage/BUS2446[13] , \iexec_stage/BUS2446[12] ,
         \iexec_stage/BUS2446[11] , \iexec_stage/BUS2446[10] ,
         \iexec_stage/BUS2446[9] , \iexec_stage/BUS2446[8] ,
         \iexec_stage/BUS2446[7] , \iexec_stage/BUS2446[6] ,
         \iexec_stage/BUS2446[5] , \iexec_stage/BUS2446[4] ,
         \iexec_stage/BUS2446[3] , \iexec_stage/BUS468[31] ,
         \iexec_stage/BUS468[15] , \iexec_stage/BUS468[9] ,
         \iexec_stage/BUS468[1] , \iexec_stage/BUS476[31] ,
         \iexec_stage/BUS476[30] , \iexec_stage/BUS476[29] ,
         \iexec_stage/BUS476[28] , \iexec_stage/BUS476[27] ,
         \iexec_stage/BUS476[26] , \iexec_stage/BUS476[25] ,
         \iexec_stage/BUS476[24] , \iexec_stage/BUS476[23] ,
         \iexec_stage/BUS476[22] , \iexec_stage/BUS476[21] ,
         \iexec_stage/BUS476[20] , \iexec_stage/BUS476[19] ,
         \iexec_stage/BUS476[18] , \iexec_stage/BUS476[17] ,
         \iexec_stage/BUS476[16] , \iexec_stage/BUS476[15] ,
         \iexec_stage/BUS476[14] , \iexec_stage/BUS476[13] ,
         \iexec_stage/BUS476[12] , \iexec_stage/BUS476[11] ,
         \iexec_stage/BUS476[10] , \iexec_stage/BUS476[9] ,
         \iexec_stage/BUS476[8] , \iexec_stage/BUS476[7] ,
         \iexec_stage/BUS476[6] , \iexec_stage/BUS476[5] ,
         \iexec_stage/BUS476[4] , \iexec_stage/BUS476[3] ,
         \iexec_stage/BUS476[2] , \iexec_stage/BUS476[1] ,
         \iexec_stage/BUS476[0] , \decoder_pipe/BUS2110[1] ,
         \decoder_pipe/BUS2110[0] , \decoder_pipe/BUS2102[2] ,
         \decoder_pipe/BUS2102[1] , \decoder_pipe/BUS2102[0] ,
         \decoder_pipe/BUS2094[1] , \decoder_pipe/BUS2094[0] ,
         \decoder_pipe/BUS2086[1] , \decoder_pipe/BUS2086[0] ,
         \decoder_pipe/BUS2072[2] , \decoder_pipe/BUS2072[0] ,
         \decoder_pipe/BUS2064[2] , \decoder_pipe/BUS2064[1] ,
         \decoder_pipe/BUS2056[2] , \decoder_pipe/BUS2056[1] ,
         \decoder_pipe/BUS2056[0] , \decoder_pipe/BUS2040[4] ,
         \decoder_pipe/BUS2040[3] , \decoder_pipe/BUS2040[2] ,
         \decoder_pipe/BUS2040[1] , \decoder_pipe/BUS2040[0] ,
         \iforward/BUS937[4] , \iforward/BUS937[3] , \iforward/BUS937[2] ,
         \iforward/BUS937[1] , \iforward/BUS937[0] , \iforward/BUS82[4] ,
         \iforward/BUS82[3] , \iforward/BUS82[2] , \iforward/BUS82[1] ,
         \iforward/BUS82[0] , \iRF_stage/MAIN_FSM/n57 ,
         \iRF_stage/MAIN_FSM/n17 , \iRF_stage/MAIN_FSM/N52 ,
         \iRF_stage/MAIN_FSM/N51 , \iRF_stage/MAIN_FSM/N50 ,
         \iRF_stage/MAIN_FSM/N37 , \iRF_stage/MAIN_FSM/N36 ,
         \iRF_stage/MAIN_FSM/N35 , \iRF_stage/MAIN_FSM/N34 ,
         \iRF_stage/MAIN_FSM/N33 , \iRF_stage/MAIN_FSM/delay_counter[0] ,
         \iRF_stage/MAIN_FSM/delay_counter[1] ,
         \iRF_stage/MAIN_FSM/delay_counter[2] ,
         \iRF_stage/MAIN_FSM/delay_counter[3] ,
         \iRF_stage/MAIN_FSM/delay_counter[4] ,
         \iRF_stage/MAIN_FSM/CurrState[0] , \iRF_stage/MAIN_FSM/CurrState[1] ,
         \iRF_stage/MAIN_FSM/CurrState[2] , \iRF_stage/i_pc_gen/N65 ,
         \iRF_stage/i_pc_gen/N64 , \iRF_stage/i_pc_gen/N63 ,
         \iRF_stage/i_pc_gen/N62 , \iRF_stage/i_pc_gen/N61 ,
         \iRF_stage/i_pc_gen/N60 , \iRF_stage/i_pc_gen/N59 ,
         \iRF_stage/i_pc_gen/N58 , \iRF_stage/i_pc_gen/N57 ,
         \iRF_stage/i_pc_gen/N56 , \iRF_stage/i_pc_gen/N55 ,
         \iRF_stage/i_pc_gen/N54 , \iRF_stage/i_pc_gen/N53 ,
         \iRF_stage/i_pc_gen/N52 , \iRF_stage/i_pc_gen/N51 ,
         \iRF_stage/i_pc_gen/N50 , \iRF_stage/i_pc_gen/N49 ,
         \iRF_stage/i_pc_gen/N48 , \iRF_stage/i_pc_gen/N47 ,
         \iRF_stage/i_pc_gen/N46 , \iRF_stage/i_pc_gen/N45 ,
         \iRF_stage/i_pc_gen/N44 , \iRF_stage/i_pc_gen/N43 ,
         \iRF_stage/i_pc_gen/N42 , \iRF_stage/i_pc_gen/N41 ,
         \iRF_stage/i_pc_gen/N40 , \iRF_stage/i_pc_gen/N39 ,
         \iRF_stage/i_pc_gen/N38 , \iRF_stage/i_pc_gen/N37 ,
         \iRF_stage/i_pc_gen/N34 , \iRF_stage/i_pc_gen/br_addr[31] ,
         \iRF_stage/i_pc_gen/br_addr[30] , \iRF_stage/i_pc_gen/br_addr[29] ,
         \iRF_stage/i_pc_gen/br_addr[28] , \iRF_stage/i_pc_gen/br_addr[27] ,
         \iRF_stage/i_pc_gen/br_addr[26] , \iRF_stage/i_pc_gen/br_addr[25] ,
         \iRF_stage/i_pc_gen/br_addr[24] , \iRF_stage/i_pc_gen/br_addr[23] ,
         \iRF_stage/i_pc_gen/br_addr[22] , \iRF_stage/i_pc_gen/br_addr[21] ,
         \iRF_stage/i_pc_gen/br_addr[20] , \iRF_stage/i_pc_gen/br_addr[19] ,
         \iRF_stage/i_pc_gen/br_addr[18] , \iRF_stage/i_pc_gen/br_addr[17] ,
         \iRF_stage/i_pc_gen/br_addr[16] , \iRF_stage/i_pc_gen/br_addr[15] ,
         \iRF_stage/i_pc_gen/br_addr[14] , \iRF_stage/i_pc_gen/br_addr[13] ,
         \iRF_stage/i_pc_gen/br_addr[12] , \iRF_stage/i_pc_gen/br_addr[11] ,
         \iRF_stage/i_pc_gen/br_addr[10] , \iRF_stage/i_pc_gen/br_addr[9] ,
         \iRF_stage/i_pc_gen/br_addr[8] , \iRF_stage/i_pc_gen/br_addr[7] ,
         \iRF_stage/i_pc_gen/br_addr[6] , \iRF_stage/i_pc_gen/br_addr[5] ,
         \iRF_stage/i_pc_gen/br_addr[4] , \iRF_stage/i_pc_gen/br_addr[3] ,
         \iRF_stage/i_pc_gen/br_addr[2] , \iRF_stage/i_pc_gen/br_addr[1] ,
         \iRF_stage/i_pc_gen/br_addr[0] , \iRF_stage/reg_bank/n1801 ,
         \iRF_stage/reg_bank/n1800 , \iRF_stage/reg_bank/n1799 ,
         \iRF_stage/reg_bank/n1798 , \iRF_stage/reg_bank/n1797 ,
         \iRF_stage/reg_bank/n1796 , \iRF_stage/reg_bank/n1795 ,
         \iRF_stage/reg_bank/n1794 , \iRF_stage/reg_bank/n1793 ,
         \iRF_stage/reg_bank/n1792 , \iRF_stage/reg_bank/n1791 ,
         \iRF_stage/reg_bank/n1790 , \iRF_stage/reg_bank/n1789 ,
         \iRF_stage/reg_bank/n1788 , \iRF_stage/reg_bank/n1787 ,
         \iRF_stage/reg_bank/n1786 , \iRF_stage/reg_bank/n1785 ,
         \iRF_stage/reg_bank/n1784 , \iRF_stage/reg_bank/n1783 ,
         \iRF_stage/reg_bank/n1782 , \iRF_stage/reg_bank/n1781 ,
         \iRF_stage/reg_bank/n1780 , \iRF_stage/reg_bank/n1779 ,
         \iRF_stage/reg_bank/n1778 , \iRF_stage/reg_bank/n1777 ,
         \iRF_stage/reg_bank/n1776 , \iRF_stage/reg_bank/n1775 ,
         \iRF_stage/reg_bank/n1774 , \iRF_stage/reg_bank/n1773 ,
         \iRF_stage/reg_bank/n1772 , \iRF_stage/reg_bank/n1771 ,
         \iRF_stage/reg_bank/n1770 , \iRF_stage/reg_bank/n1769 ,
         \iRF_stage/reg_bank/n1768 , \iRF_stage/reg_bank/n1767 ,
         \iRF_stage/reg_bank/n1766 , \iRF_stage/reg_bank/n1765 ,
         \iRF_stage/reg_bank/n1764 , \iRF_stage/reg_bank/n1763 ,
         \iRF_stage/reg_bank/n1762 , \iRF_stage/reg_bank/n1761 ,
         \iRF_stage/reg_bank/n1760 , \iRF_stage/reg_bank/n1759 ,
         \iRF_stage/reg_bank/n1758 , \iRF_stage/reg_bank/n1757 ,
         \iRF_stage/reg_bank/n1756 , \iRF_stage/reg_bank/n1755 ,
         \iRF_stage/reg_bank/n1754 , \iRF_stage/reg_bank/n1753 ,
         \iRF_stage/reg_bank/n1752 , \iRF_stage/reg_bank/n1751 ,
         \iRF_stage/reg_bank/n1750 , \iRF_stage/reg_bank/n1749 ,
         \iRF_stage/reg_bank/n1748 , \iRF_stage/reg_bank/n1747 ,
         \iRF_stage/reg_bank/n1746 , \iRF_stage/reg_bank/n1745 ,
         \iRF_stage/reg_bank/n1744 , \iRF_stage/reg_bank/n1743 ,
         \iRF_stage/reg_bank/n1742 , \iRF_stage/reg_bank/n1741 ,
         \iRF_stage/reg_bank/n1740 , \iRF_stage/reg_bank/n1739 ,
         \iRF_stage/reg_bank/n1738 , \iRF_stage/reg_bank/n1737 ,
         \iRF_stage/reg_bank/n1736 , \iRF_stage/reg_bank/n1735 ,
         \iRF_stage/reg_bank/n1734 , \iRF_stage/reg_bank/n1733 ,
         \iRF_stage/reg_bank/n1732 , \iRF_stage/reg_bank/n1731 ,
         \iRF_stage/reg_bank/n1730 , \iRF_stage/reg_bank/n1729 ,
         \iRF_stage/reg_bank/n1728 , \iRF_stage/reg_bank/n1727 ,
         \iRF_stage/reg_bank/n1726 , \iRF_stage/reg_bank/n1725 ,
         \iRF_stage/reg_bank/n1724 , \iRF_stage/reg_bank/n1723 ,
         \iRF_stage/reg_bank/n1722 , \iRF_stage/reg_bank/n1721 ,
         \iRF_stage/reg_bank/n1720 , \iRF_stage/reg_bank/n1719 ,
         \iRF_stage/reg_bank/n1718 , \iRF_stage/reg_bank/n1717 ,
         \iRF_stage/reg_bank/n1716 , \iRF_stage/reg_bank/n1715 ,
         \iRF_stage/reg_bank/n1714 , \iRF_stage/reg_bank/n1713 ,
         \iRF_stage/reg_bank/n1712 , \iRF_stage/reg_bank/n1711 ,
         \iRF_stage/reg_bank/n1710 , \iRF_stage/reg_bank/n1709 ,
         \iRF_stage/reg_bank/n1708 , \iRF_stage/reg_bank/n1707 ,
         \iRF_stage/reg_bank/n1706 , \iRF_stage/reg_bank/n1705 ,
         \iRF_stage/reg_bank/n1704 , \iRF_stage/reg_bank/n1703 ,
         \iRF_stage/reg_bank/n1702 , \iRF_stage/reg_bank/n1701 ,
         \iRF_stage/reg_bank/n1700 , \iRF_stage/reg_bank/n1699 ,
         \iRF_stage/reg_bank/n1698 , \iRF_stage/reg_bank/n1697 ,
         \iRF_stage/reg_bank/n1696 , \iRF_stage/reg_bank/n1695 ,
         \iRF_stage/reg_bank/n1694 , \iRF_stage/reg_bank/n1693 ,
         \iRF_stage/reg_bank/n1692 , \iRF_stage/reg_bank/n1691 ,
         \iRF_stage/reg_bank/n1690 , \iRF_stage/reg_bank/n1689 ,
         \iRF_stage/reg_bank/n1688 , \iRF_stage/reg_bank/n1687 ,
         \iRF_stage/reg_bank/n1686 , \iRF_stage/reg_bank/n1685 ,
         \iRF_stage/reg_bank/n1684 , \iRF_stage/reg_bank/n1683 ,
         \iRF_stage/reg_bank/n1682 , \iRF_stage/reg_bank/n1681 ,
         \iRF_stage/reg_bank/n1680 , \iRF_stage/reg_bank/n1679 ,
         \iRF_stage/reg_bank/n1678 , \iRF_stage/reg_bank/n1677 ,
         \iRF_stage/reg_bank/n1676 , \iRF_stage/reg_bank/n1675 ,
         \iRF_stage/reg_bank/n1674 , \iRF_stage/reg_bank/n1673 ,
         \iRF_stage/reg_bank/n1672 , \iRF_stage/reg_bank/n1671 ,
         \iRF_stage/reg_bank/n1670 , \iRF_stage/reg_bank/n1669 ,
         \iRF_stage/reg_bank/n1668 , \iRF_stage/reg_bank/n1667 ,
         \iRF_stage/reg_bank/n1666 , \iRF_stage/reg_bank/n1665 ,
         \iRF_stage/reg_bank/n1664 , \iRF_stage/reg_bank/n1663 ,
         \iRF_stage/reg_bank/n1662 , \iRF_stage/reg_bank/n1661 ,
         \iRF_stage/reg_bank/n1660 , \iRF_stage/reg_bank/n1659 ,
         \iRF_stage/reg_bank/n1658 , \iRF_stage/reg_bank/n1657 ,
         \iRF_stage/reg_bank/n1656 , \iRF_stage/reg_bank/n1655 ,
         \iRF_stage/reg_bank/n1654 , \iRF_stage/reg_bank/n1653 ,
         \iRF_stage/reg_bank/n1652 , \iRF_stage/reg_bank/n1651 ,
         \iRF_stage/reg_bank/n1650 , \iRF_stage/reg_bank/n1649 ,
         \iRF_stage/reg_bank/n1648 , \iRF_stage/reg_bank/n1647 ,
         \iRF_stage/reg_bank/n1646 , \iRF_stage/reg_bank/n1645 ,
         \iRF_stage/reg_bank/n1644 , \iRF_stage/reg_bank/n1643 ,
         \iRF_stage/reg_bank/n1642 , \iRF_stage/reg_bank/n1641 ,
         \iRF_stage/reg_bank/n1640 , \iRF_stage/reg_bank/n1639 ,
         \iRF_stage/reg_bank/n1638 , \iRF_stage/reg_bank/n1637 ,
         \iRF_stage/reg_bank/n1636 , \iRF_stage/reg_bank/n1635 ,
         \iRF_stage/reg_bank/n1634 , \iRF_stage/reg_bank/n1633 ,
         \iRF_stage/reg_bank/n1632 , \iRF_stage/reg_bank/n1631 ,
         \iRF_stage/reg_bank/n1630 , \iRF_stage/reg_bank/n1629 ,
         \iRF_stage/reg_bank/n1628 , \iRF_stage/reg_bank/n1627 ,
         \iRF_stage/reg_bank/n1626 , \iRF_stage/reg_bank/n1625 ,
         \iRF_stage/reg_bank/n1624 , \iRF_stage/reg_bank/n1623 ,
         \iRF_stage/reg_bank/n1622 , \iRF_stage/reg_bank/n1621 ,
         \iRF_stage/reg_bank/n1620 , \iRF_stage/reg_bank/n1619 ,
         \iRF_stage/reg_bank/n1618 , \iRF_stage/reg_bank/n1617 ,
         \iRF_stage/reg_bank/n1616 , \iRF_stage/reg_bank/n1615 ,
         \iRF_stage/reg_bank/n1614 , \iRF_stage/reg_bank/n1613 ,
         \iRF_stage/reg_bank/n1612 , \iRF_stage/reg_bank/n1611 ,
         \iRF_stage/reg_bank/n1610 , \iRF_stage/reg_bank/n1609 ,
         \iRF_stage/reg_bank/n1608 , \iRF_stage/reg_bank/n1607 ,
         \iRF_stage/reg_bank/n1606 , \iRF_stage/reg_bank/n1605 ,
         \iRF_stage/reg_bank/n1604 , \iRF_stage/reg_bank/n1603 ,
         \iRF_stage/reg_bank/n1602 , \iRF_stage/reg_bank/n1601 ,
         \iRF_stage/reg_bank/n1600 , \iRF_stage/reg_bank/n1599 ,
         \iRF_stage/reg_bank/n1598 , \iRF_stage/reg_bank/n1597 ,
         \iRF_stage/reg_bank/n1596 , \iRF_stage/reg_bank/n1595 ,
         \iRF_stage/reg_bank/n1594 , \iRF_stage/reg_bank/n1593 ,
         \iRF_stage/reg_bank/n1592 , \iRF_stage/reg_bank/n1591 ,
         \iRF_stage/reg_bank/n1590 , \iRF_stage/reg_bank/n1589 ,
         \iRF_stage/reg_bank/n1588 , \iRF_stage/reg_bank/n1587 ,
         \iRF_stage/reg_bank/n1586 , \iRF_stage/reg_bank/n1585 ,
         \iRF_stage/reg_bank/n1584 , \iRF_stage/reg_bank/n1583 ,
         \iRF_stage/reg_bank/n1582 , \iRF_stage/reg_bank/n1581 ,
         \iRF_stage/reg_bank/n1580 , \iRF_stage/reg_bank/n1579 ,
         \iRF_stage/reg_bank/n1578 , \iRF_stage/reg_bank/n1577 ,
         \iRF_stage/reg_bank/n1576 , \iRF_stage/reg_bank/n1575 ,
         \iRF_stage/reg_bank/n1574 , \iRF_stage/reg_bank/n1573 ,
         \iRF_stage/reg_bank/n1572 , \iRF_stage/reg_bank/n1571 ,
         \iRF_stage/reg_bank/n1570 , \iRF_stage/reg_bank/n1569 ,
         \iRF_stage/reg_bank/n1568 , \iRF_stage/reg_bank/n1567 ,
         \iRF_stage/reg_bank/n1566 , \iRF_stage/reg_bank/n1565 ,
         \iRF_stage/reg_bank/n1564 , \iRF_stage/reg_bank/n1563 ,
         \iRF_stage/reg_bank/n1562 , \iRF_stage/reg_bank/n1561 ,
         \iRF_stage/reg_bank/n1560 , \iRF_stage/reg_bank/n1559 ,
         \iRF_stage/reg_bank/n1558 , \iRF_stage/reg_bank/n1557 ,
         \iRF_stage/reg_bank/n1556 , \iRF_stage/reg_bank/n1555 ,
         \iRF_stage/reg_bank/n1554 , \iRF_stage/reg_bank/n1553 ,
         \iRF_stage/reg_bank/n1552 , \iRF_stage/reg_bank/n1551 ,
         \iRF_stage/reg_bank/n1550 , \iRF_stage/reg_bank/n1549 ,
         \iRF_stage/reg_bank/n1548 , \iRF_stage/reg_bank/n1547 ,
         \iRF_stage/reg_bank/n1546 , \iRF_stage/reg_bank/n1545 ,
         \iRF_stage/reg_bank/n1544 , \iRF_stage/reg_bank/n1543 ,
         \iRF_stage/reg_bank/n1542 , \iRF_stage/reg_bank/n1541 ,
         \iRF_stage/reg_bank/n1540 , \iRF_stage/reg_bank/n1539 ,
         \iRF_stage/reg_bank/n1538 , \iRF_stage/reg_bank/n1537 ,
         \iRF_stage/reg_bank/n1536 , \iRF_stage/reg_bank/n1535 ,
         \iRF_stage/reg_bank/n1534 , \iRF_stage/reg_bank/n1533 ,
         \iRF_stage/reg_bank/n1532 , \iRF_stage/reg_bank/n1531 ,
         \iRF_stage/reg_bank/n1530 , \iRF_stage/reg_bank/n1529 ,
         \iRF_stage/reg_bank/n1528 , \iRF_stage/reg_bank/n1527 ,
         \iRF_stage/reg_bank/n1526 , \iRF_stage/reg_bank/n1525 ,
         \iRF_stage/reg_bank/n1524 , \iRF_stage/reg_bank/n1523 ,
         \iRF_stage/reg_bank/n1522 , \iRF_stage/reg_bank/n1521 ,
         \iRF_stage/reg_bank/n1520 , \iRF_stage/reg_bank/n1519 ,
         \iRF_stage/reg_bank/n1518 , \iRF_stage/reg_bank/n1517 ,
         \iRF_stage/reg_bank/n1516 , \iRF_stage/reg_bank/n1515 ,
         \iRF_stage/reg_bank/n1514 , \iRF_stage/reg_bank/n1513 ,
         \iRF_stage/reg_bank/n1512 , \iRF_stage/reg_bank/n1511 ,
         \iRF_stage/reg_bank/n1510 , \iRF_stage/reg_bank/n1509 ,
         \iRF_stage/reg_bank/n1508 , \iRF_stage/reg_bank/n1507 ,
         \iRF_stage/reg_bank/n1506 , \iRF_stage/reg_bank/n1505 ,
         \iRF_stage/reg_bank/n1504 , \iRF_stage/reg_bank/n1503 ,
         \iRF_stage/reg_bank/n1502 , \iRF_stage/reg_bank/n1501 ,
         \iRF_stage/reg_bank/n1500 , \iRF_stage/reg_bank/n1499 ,
         \iRF_stage/reg_bank/n1498 , \iRF_stage/reg_bank/n1497 ,
         \iRF_stage/reg_bank/n1496 , \iRF_stage/reg_bank/n1495 ,
         \iRF_stage/reg_bank/n1494 , \iRF_stage/reg_bank/n1493 ,
         \iRF_stage/reg_bank/n1492 , \iRF_stage/reg_bank/n1491 ,
         \iRF_stage/reg_bank/n1490 , \iRF_stage/reg_bank/n1489 ,
         \iRF_stage/reg_bank/n1488 , \iRF_stage/reg_bank/n1487 ,
         \iRF_stage/reg_bank/n1486 , \iRF_stage/reg_bank/n1485 ,
         \iRF_stage/reg_bank/n1484 , \iRF_stage/reg_bank/n1483 ,
         \iRF_stage/reg_bank/n1482 , \iRF_stage/reg_bank/n1481 ,
         \iRF_stage/reg_bank/n1480 , \iRF_stage/reg_bank/n1479 ,
         \iRF_stage/reg_bank/n1478 , \iRF_stage/reg_bank/n1477 ,
         \iRF_stage/reg_bank/n1476 , \iRF_stage/reg_bank/n1475 ,
         \iRF_stage/reg_bank/n1474 , \iRF_stage/reg_bank/n1473 ,
         \iRF_stage/reg_bank/n1472 , \iRF_stage/reg_bank/n1471 ,
         \iRF_stage/reg_bank/n1470 , \iRF_stage/reg_bank/n1469 ,
         \iRF_stage/reg_bank/n1468 , \iRF_stage/reg_bank/n1467 ,
         \iRF_stage/reg_bank/n1466 , \iRF_stage/reg_bank/n1465 ,
         \iRF_stage/reg_bank/n1464 , \iRF_stage/reg_bank/n1463 ,
         \iRF_stage/reg_bank/n1462 , \iRF_stage/reg_bank/n1461 ,
         \iRF_stage/reg_bank/n1460 , \iRF_stage/reg_bank/n1459 ,
         \iRF_stage/reg_bank/n1458 , \iRF_stage/reg_bank/n1457 ,
         \iRF_stage/reg_bank/n1456 , \iRF_stage/reg_bank/n1455 ,
         \iRF_stage/reg_bank/n1454 , \iRF_stage/reg_bank/n1453 ,
         \iRF_stage/reg_bank/n1452 , \iRF_stage/reg_bank/n1451 ,
         \iRF_stage/reg_bank/n1450 , \iRF_stage/reg_bank/n1449 ,
         \iRF_stage/reg_bank/n1448 , \iRF_stage/reg_bank/n1447 ,
         \iRF_stage/reg_bank/n1446 , \iRF_stage/reg_bank/n1445 ,
         \iRF_stage/reg_bank/n1444 , \iRF_stage/reg_bank/n1443 ,
         \iRF_stage/reg_bank/n1442 , \iRF_stage/reg_bank/n1441 ,
         \iRF_stage/reg_bank/n1440 , \iRF_stage/reg_bank/n1439 ,
         \iRF_stage/reg_bank/n1438 , \iRF_stage/reg_bank/n1437 ,
         \iRF_stage/reg_bank/n1436 , \iRF_stage/reg_bank/n1435 ,
         \iRF_stage/reg_bank/n1434 , \iRF_stage/reg_bank/n1433 ,
         \iRF_stage/reg_bank/n1432 , \iRF_stage/reg_bank/n1431 ,
         \iRF_stage/reg_bank/n1430 , \iRF_stage/reg_bank/n1429 ,
         \iRF_stage/reg_bank/n1428 , \iRF_stage/reg_bank/n1427 ,
         \iRF_stage/reg_bank/n1426 , \iRF_stage/reg_bank/n1425 ,
         \iRF_stage/reg_bank/n1424 , \iRF_stage/reg_bank/n1423 ,
         \iRF_stage/reg_bank/n1422 , \iRF_stage/reg_bank/n1421 ,
         \iRF_stage/reg_bank/n1420 , \iRF_stage/reg_bank/n1419 ,
         \iRF_stage/reg_bank/n1418 , \iRF_stage/reg_bank/n1417 ,
         \iRF_stage/reg_bank/n1416 , \iRF_stage/reg_bank/n1415 ,
         \iRF_stage/reg_bank/n1414 , \iRF_stage/reg_bank/n1413 ,
         \iRF_stage/reg_bank/n1412 , \iRF_stage/reg_bank/n1411 ,
         \iRF_stage/reg_bank/n1410 , \iRF_stage/reg_bank/n1409 ,
         \iRF_stage/reg_bank/n1408 , \iRF_stage/reg_bank/n1407 ,
         \iRF_stage/reg_bank/n1406 , \iRF_stage/reg_bank/n1405 ,
         \iRF_stage/reg_bank/n1404 , \iRF_stage/reg_bank/n1403 ,
         \iRF_stage/reg_bank/n1402 , \iRF_stage/reg_bank/n1401 ,
         \iRF_stage/reg_bank/n1400 , \iRF_stage/reg_bank/n1399 ,
         \iRF_stage/reg_bank/n1398 , \iRF_stage/reg_bank/n1397 ,
         \iRF_stage/reg_bank/n1396 , \iRF_stage/reg_bank/n1395 ,
         \iRF_stage/reg_bank/n1394 , \iRF_stage/reg_bank/n1393 ,
         \iRF_stage/reg_bank/n1392 , \iRF_stage/reg_bank/n1391 ,
         \iRF_stage/reg_bank/n1390 , \iRF_stage/reg_bank/n1389 ,
         \iRF_stage/reg_bank/n1388 , \iRF_stage/reg_bank/n1387 ,
         \iRF_stage/reg_bank/n1386 , \iRF_stage/reg_bank/n1385 ,
         \iRF_stage/reg_bank/n1384 , \iRF_stage/reg_bank/n1383 ,
         \iRF_stage/reg_bank/n1382 , \iRF_stage/reg_bank/n1381 ,
         \iRF_stage/reg_bank/n1380 , \iRF_stage/reg_bank/n1379 ,
         \iRF_stage/reg_bank/n1378 , \iRF_stage/reg_bank/n1377 ,
         \iRF_stage/reg_bank/n1376 , \iRF_stage/reg_bank/n1375 ,
         \iRF_stage/reg_bank/n1374 , \iRF_stage/reg_bank/n1373 ,
         \iRF_stage/reg_bank/n1372 , \iRF_stage/reg_bank/n1371 ,
         \iRF_stage/reg_bank/n1370 , \iRF_stage/reg_bank/n1369 ,
         \iRF_stage/reg_bank/n1368 , \iRF_stage/reg_bank/n1367 ,
         \iRF_stage/reg_bank/n1366 , \iRF_stage/reg_bank/n1365 ,
         \iRF_stage/reg_bank/n1364 , \iRF_stage/reg_bank/n1363 ,
         \iRF_stage/reg_bank/n1362 , \iRF_stage/reg_bank/n1361 ,
         \iRF_stage/reg_bank/n1360 , \iRF_stage/reg_bank/n1359 ,
         \iRF_stage/reg_bank/n1358 , \iRF_stage/reg_bank/n1357 ,
         \iRF_stage/reg_bank/n1356 , \iRF_stage/reg_bank/n1355 ,
         \iRF_stage/reg_bank/n1354 , \iRF_stage/reg_bank/n1353 ,
         \iRF_stage/reg_bank/n1352 , \iRF_stage/reg_bank/n1351 ,
         \iRF_stage/reg_bank/n1350 , \iRF_stage/reg_bank/n1349 ,
         \iRF_stage/reg_bank/n1348 , \iRF_stage/reg_bank/n1347 ,
         \iRF_stage/reg_bank/n1346 , \iRF_stage/reg_bank/n1345 ,
         \iRF_stage/reg_bank/n1344 , \iRF_stage/reg_bank/n1343 ,
         \iRF_stage/reg_bank/n1342 , \iRF_stage/reg_bank/n1341 ,
         \iRF_stage/reg_bank/n1340 , \iRF_stage/reg_bank/n1339 ,
         \iRF_stage/reg_bank/n1338 , \iRF_stage/reg_bank/n1337 ,
         \iRF_stage/reg_bank/n1336 , \iRF_stage/reg_bank/n1335 ,
         \iRF_stage/reg_bank/n1334 , \iRF_stage/reg_bank/n1333 ,
         \iRF_stage/reg_bank/n1332 , \iRF_stage/reg_bank/n1331 ,
         \iRF_stage/reg_bank/n1330 , \iRF_stage/reg_bank/n1329 ,
         \iRF_stage/reg_bank/n1328 , \iRF_stage/reg_bank/n1327 ,
         \iRF_stage/reg_bank/n1326 , \iRF_stage/reg_bank/n1325 ,
         \iRF_stage/reg_bank/n1324 , \iRF_stage/reg_bank/n1323 ,
         \iRF_stage/reg_bank/n1322 , \iRF_stage/reg_bank/n1321 ,
         \iRF_stage/reg_bank/n1320 , \iRF_stage/reg_bank/n1319 ,
         \iRF_stage/reg_bank/n1318 , \iRF_stage/reg_bank/n1317 ,
         \iRF_stage/reg_bank/n1316 , \iRF_stage/reg_bank/n1315 ,
         \iRF_stage/reg_bank/n1314 , \iRF_stage/reg_bank/n1313 ,
         \iRF_stage/reg_bank/n1312 , \iRF_stage/reg_bank/n1311 ,
         \iRF_stage/reg_bank/n1310 , \iRF_stage/reg_bank/n1309 ,
         \iRF_stage/reg_bank/n1308 , \iRF_stage/reg_bank/n1307 ,
         \iRF_stage/reg_bank/n1306 , \iRF_stage/reg_bank/n1305 ,
         \iRF_stage/reg_bank/n1304 , \iRF_stage/reg_bank/n1303 ,
         \iRF_stage/reg_bank/n1302 , \iRF_stage/reg_bank/n1301 ,
         \iRF_stage/reg_bank/n1300 , \iRF_stage/reg_bank/n1299 ,
         \iRF_stage/reg_bank/n1298 , \iRF_stage/reg_bank/n1297 ,
         \iRF_stage/reg_bank/n1296 , \iRF_stage/reg_bank/n1295 ,
         \iRF_stage/reg_bank/n1294 , \iRF_stage/reg_bank/n1293 ,
         \iRF_stage/reg_bank/n1292 , \iRF_stage/reg_bank/n1291 ,
         \iRF_stage/reg_bank/n1290 , \iRF_stage/reg_bank/n1289 ,
         \iRF_stage/reg_bank/n1288 , \iRF_stage/reg_bank/n1287 ,
         \iRF_stage/reg_bank/n1286 , \iRF_stage/reg_bank/n1285 ,
         \iRF_stage/reg_bank/n1284 , \iRF_stage/reg_bank/n1283 ,
         \iRF_stage/reg_bank/n1282 , \iRF_stage/reg_bank/n1281 ,
         \iRF_stage/reg_bank/n1280 , \iRF_stage/reg_bank/n1279 ,
         \iRF_stage/reg_bank/n1278 , \iRF_stage/reg_bank/n1277 ,
         \iRF_stage/reg_bank/n1276 , \iRF_stage/reg_bank/n1275 ,
         \iRF_stage/reg_bank/n1274 , \iRF_stage/reg_bank/n1273 ,
         \iRF_stage/reg_bank/n1272 , \iRF_stage/reg_bank/n1271 ,
         \iRF_stage/reg_bank/n1270 , \iRF_stage/reg_bank/n1269 ,
         \iRF_stage/reg_bank/n1268 , \iRF_stage/reg_bank/n1267 ,
         \iRF_stage/reg_bank/n1266 , \iRF_stage/reg_bank/n1265 ,
         \iRF_stage/reg_bank/n1264 , \iRF_stage/reg_bank/n1263 ,
         \iRF_stage/reg_bank/n1262 , \iRF_stage/reg_bank/n1261 ,
         \iRF_stage/reg_bank/n1260 , \iRF_stage/reg_bank/n1259 ,
         \iRF_stage/reg_bank/n1258 , \iRF_stage/reg_bank/n1257 ,
         \iRF_stage/reg_bank/n1256 , \iRF_stage/reg_bank/n1255 ,
         \iRF_stage/reg_bank/n1254 , \iRF_stage/reg_bank/n1253 ,
         \iRF_stage/reg_bank/n1252 , \iRF_stage/reg_bank/n1251 ,
         \iRF_stage/reg_bank/n1250 , \iRF_stage/reg_bank/n1249 ,
         \iRF_stage/reg_bank/n1248 , \iRF_stage/reg_bank/n1247 ,
         \iRF_stage/reg_bank/n1246 , \iRF_stage/reg_bank/n1245 ,
         \iRF_stage/reg_bank/n1244 , \iRF_stage/reg_bank/n1243 ,
         \iRF_stage/reg_bank/n1242 , \iRF_stage/reg_bank/n1241 ,
         \iRF_stage/reg_bank/n1240 , \iRF_stage/reg_bank/n1239 ,
         \iRF_stage/reg_bank/n1238 , \iRF_stage/reg_bank/n1237 ,
         \iRF_stage/reg_bank/n1236 , \iRF_stage/reg_bank/n1235 ,
         \iRF_stage/reg_bank/n1234 , \iRF_stage/reg_bank/n1233 ,
         \iRF_stage/reg_bank/n1232 , \iRF_stage/reg_bank/n1231 ,
         \iRF_stage/reg_bank/n1230 , \iRF_stage/reg_bank/n1229 ,
         \iRF_stage/reg_bank/n1228 , \iRF_stage/reg_bank/n1227 ,
         \iRF_stage/reg_bank/n1226 , \iRF_stage/reg_bank/n1225 ,
         \iRF_stage/reg_bank/n1224 , \iRF_stage/reg_bank/n1223 ,
         \iRF_stage/reg_bank/n1222 , \iRF_stage/reg_bank/n1221 ,
         \iRF_stage/reg_bank/n1220 , \iRF_stage/reg_bank/n1219 ,
         \iRF_stage/reg_bank/n1218 , \iRF_stage/reg_bank/n1217 ,
         \iRF_stage/reg_bank/n1216 , \iRF_stage/reg_bank/n1215 ,
         \iRF_stage/reg_bank/n1214 , \iRF_stage/reg_bank/n1213 ,
         \iRF_stage/reg_bank/n1212 , \iRF_stage/reg_bank/n1211 ,
         \iRF_stage/reg_bank/n1210 , \iRF_stage/reg_bank/n1209 ,
         \iRF_stage/reg_bank/n1208 , \iRF_stage/reg_bank/n1207 ,
         \iRF_stage/reg_bank/n1206 , \iRF_stage/reg_bank/n1205 ,
         \iRF_stage/reg_bank/n1204 , \iRF_stage/reg_bank/n1203 ,
         \iRF_stage/reg_bank/n1202 , \iRF_stage/reg_bank/n1201 ,
         \iRF_stage/reg_bank/n1200 , \iRF_stage/reg_bank/n1199 ,
         \iRF_stage/reg_bank/n1198 , \iRF_stage/reg_bank/n1197 ,
         \iRF_stage/reg_bank/n1196 , \iRF_stage/reg_bank/n1195 ,
         \iRF_stage/reg_bank/n1194 , \iRF_stage/reg_bank/n1193 ,
         \iRF_stage/reg_bank/n1192 , \iRF_stage/reg_bank/n1191 ,
         \iRF_stage/reg_bank/n1190 , \iRF_stage/reg_bank/n1189 ,
         \iRF_stage/reg_bank/n1188 , \iRF_stage/reg_bank/n1187 ,
         \iRF_stage/reg_bank/n1186 , \iRF_stage/reg_bank/n1185 ,
         \iRF_stage/reg_bank/n1184 , \iRF_stage/reg_bank/n1183 ,
         \iRF_stage/reg_bank/n1182 , \iRF_stage/reg_bank/n1181 ,
         \iRF_stage/reg_bank/n1180 , \iRF_stage/reg_bank/n1179 ,
         \iRF_stage/reg_bank/n1178 , \iRF_stage/reg_bank/n1177 ,
         \iRF_stage/reg_bank/n1176 , \iRF_stage/reg_bank/n1175 ,
         \iRF_stage/reg_bank/n1174 , \iRF_stage/reg_bank/n1173 ,
         \iRF_stage/reg_bank/n1172 , \iRF_stage/reg_bank/n1171 ,
         \iRF_stage/reg_bank/n1170 , \iRF_stage/reg_bank/n1169 ,
         \iRF_stage/reg_bank/n1168 , \iRF_stage/reg_bank/n1167 ,
         \iRF_stage/reg_bank/n1166 , \iRF_stage/reg_bank/n1165 ,
         \iRF_stage/reg_bank/n1164 , \iRF_stage/reg_bank/n1163 ,
         \iRF_stage/reg_bank/n1162 , \iRF_stage/reg_bank/n1161 ,
         \iRF_stage/reg_bank/n1160 , \iRF_stage/reg_bank/n1159 ,
         \iRF_stage/reg_bank/n1158 , \iRF_stage/reg_bank/n1157 ,
         \iRF_stage/reg_bank/n1156 , \iRF_stage/reg_bank/n1155 ,
         \iRF_stage/reg_bank/n1154 , \iRF_stage/reg_bank/n1153 ,
         \iRF_stage/reg_bank/n1152 , \iRF_stage/reg_bank/n1151 ,
         \iRF_stage/reg_bank/n1150 , \iRF_stage/reg_bank/n1149 ,
         \iRF_stage/reg_bank/n1148 , \iRF_stage/reg_bank/n1147 ,
         \iRF_stage/reg_bank/n1146 , \iRF_stage/reg_bank/n1145 ,
         \iRF_stage/reg_bank/n1144 , \iRF_stage/reg_bank/n1143 ,
         \iRF_stage/reg_bank/n1142 , \iRF_stage/reg_bank/n1141 ,
         \iRF_stage/reg_bank/n1140 , \iRF_stage/reg_bank/n1139 ,
         \iRF_stage/reg_bank/n1138 , \iRF_stage/reg_bank/n1137 ,
         \iRF_stage/reg_bank/n1136 , \iRF_stage/reg_bank/n1135 ,
         \iRF_stage/reg_bank/n1134 , \iRF_stage/reg_bank/n1133 ,
         \iRF_stage/reg_bank/n1132 , \iRF_stage/reg_bank/n1131 ,
         \iRF_stage/reg_bank/n1130 , \iRF_stage/reg_bank/n1129 ,
         \iRF_stage/reg_bank/n1128 , \iRF_stage/reg_bank/n1127 ,
         \iRF_stage/reg_bank/n1126 , \iRF_stage/reg_bank/n1125 ,
         \iRF_stage/reg_bank/n1124 , \iRF_stage/reg_bank/n1123 ,
         \iRF_stage/reg_bank/n1122 , \iRF_stage/reg_bank/n1121 ,
         \iRF_stage/reg_bank/n1120 , \iRF_stage/reg_bank/n1119 ,
         \iRF_stage/reg_bank/n1118 , \iRF_stage/reg_bank/n1117 ,
         \iRF_stage/reg_bank/n1116 , \iRF_stage/reg_bank/n1115 ,
         \iRF_stage/reg_bank/n1114 , \iRF_stage/reg_bank/n1113 ,
         \iRF_stage/reg_bank/n1112 , \iRF_stage/reg_bank/n1111 ,
         \iRF_stage/reg_bank/n1110 , \iRF_stage/reg_bank/n1109 ,
         \iRF_stage/reg_bank/n1108 , \iRF_stage/reg_bank/n1107 ,
         \iRF_stage/reg_bank/n1106 , \iRF_stage/reg_bank/n1105 ,
         \iRF_stage/reg_bank/n1104 , \iRF_stage/reg_bank/n1103 ,
         \iRF_stage/reg_bank/n1102 , \iRF_stage/reg_bank/n1101 ,
         \iRF_stage/reg_bank/n1100 , \iRF_stage/reg_bank/n1099 ,
         \iRF_stage/reg_bank/n1098 , \iRF_stage/reg_bank/n1097 ,
         \iRF_stage/reg_bank/n1096 , \iRF_stage/reg_bank/n1095 ,
         \iRF_stage/reg_bank/n1094 , \iRF_stage/reg_bank/n1093 ,
         \iRF_stage/reg_bank/n1092 , \iRF_stage/reg_bank/n1091 ,
         \iRF_stage/reg_bank/n1090 , \iRF_stage/reg_bank/n1089 ,
         \iRF_stage/reg_bank/n1088 , \iRF_stage/reg_bank/n1087 ,
         \iRF_stage/reg_bank/n1086 , \iRF_stage/reg_bank/n1085 ,
         \iRF_stage/reg_bank/n1084 , \iRF_stage/reg_bank/n1083 ,
         \iRF_stage/reg_bank/n1082 , \iRF_stage/reg_bank/n1081 ,
         \iRF_stage/reg_bank/n1080 , \iRF_stage/reg_bank/n1079 ,
         \iRF_stage/reg_bank/n1078 , \iRF_stage/reg_bank/n1077 ,
         \iRF_stage/reg_bank/n1076 , \iRF_stage/reg_bank/n1075 ,
         \iRF_stage/reg_bank/n1074 , \iRF_stage/reg_bank/n1073 ,
         \iRF_stage/reg_bank/n1072 , \iRF_stage/reg_bank/n1071 ,
         \iRF_stage/reg_bank/n1070 , \iRF_stage/reg_bank/n1069 ,
         \iRF_stage/reg_bank/n1068 , \iRF_stage/reg_bank/n1067 ,
         \iRF_stage/reg_bank/n1066 , \iRF_stage/reg_bank/n1065 ,
         \iRF_stage/reg_bank/n1064 , \iRF_stage/reg_bank/n1063 ,
         \iRF_stage/reg_bank/n1062 , \iRF_stage/reg_bank/n1061 ,
         \iRF_stage/reg_bank/n1060 , \iRF_stage/reg_bank/n1059 ,
         \iRF_stage/reg_bank/n1058 , \iRF_stage/reg_bank/n1057 ,
         \iRF_stage/reg_bank/n1056 , \iRF_stage/reg_bank/n1055 ,
         \iRF_stage/reg_bank/n1054 , \iRF_stage/reg_bank/n1053 ,
         \iRF_stage/reg_bank/n1052 , \iRF_stage/reg_bank/n1051 ,
         \iRF_stage/reg_bank/n1050 , \iRF_stage/reg_bank/n1049 ,
         \iRF_stage/reg_bank/n1048 , \iRF_stage/reg_bank/n1047 ,
         \iRF_stage/reg_bank/n1046 , \iRF_stage/reg_bank/n1045 ,
         \iRF_stage/reg_bank/n1044 , \iRF_stage/reg_bank/n1043 ,
         \iRF_stage/reg_bank/n1042 , \iRF_stage/reg_bank/n1041 ,
         \iRF_stage/reg_bank/n1040 , \iRF_stage/reg_bank/n1039 ,
         \iRF_stage/reg_bank/n1038 , \iRF_stage/reg_bank/n1037 ,
         \iRF_stage/reg_bank/n1036 , \iRF_stage/reg_bank/n1035 ,
         \iRF_stage/reg_bank/n1034 , \iRF_stage/reg_bank/n1033 ,
         \iRF_stage/reg_bank/n1032 , \iRF_stage/reg_bank/n1031 ,
         \iRF_stage/reg_bank/n1030 , \iRF_stage/reg_bank/n1029 ,
         \iRF_stage/reg_bank/n1028 , \iRF_stage/reg_bank/n1027 ,
         \iRF_stage/reg_bank/n1026 , \iRF_stage/reg_bank/n1025 ,
         \iRF_stage/reg_bank/n1024 , \iRF_stage/reg_bank/n1023 ,
         \iRF_stage/reg_bank/n1022 , \iRF_stage/reg_bank/n1021 ,
         \iRF_stage/reg_bank/n1020 , \iRF_stage/reg_bank/n1019 ,
         \iRF_stage/reg_bank/n1018 , \iRF_stage/reg_bank/n1017 ,
         \iRF_stage/reg_bank/n1016 , \iRF_stage/reg_bank/n1015 ,
         \iRF_stage/reg_bank/n1014 , \iRF_stage/reg_bank/n1013 ,
         \iRF_stage/reg_bank/n1012 , \iRF_stage/reg_bank/n1011 ,
         \iRF_stage/reg_bank/n1010 , \iRF_stage/reg_bank/n1009 ,
         \iRF_stage/reg_bank/n1008 , \iRF_stage/reg_bank/n1007 ,
         \iRF_stage/reg_bank/n1006 , \iRF_stage/reg_bank/n1005 ,
         \iRF_stage/reg_bank/n1004 , \iRF_stage/reg_bank/n1003 ,
         \iRF_stage/reg_bank/n1002 , \iRF_stage/reg_bank/n1001 ,
         \iRF_stage/reg_bank/n1000 , \iRF_stage/reg_bank/n999 ,
         \iRF_stage/reg_bank/n998 , \iRF_stage/reg_bank/n997 ,
         \iRF_stage/reg_bank/n996 , \iRF_stage/reg_bank/n995 ,
         \iRF_stage/reg_bank/n994 , \iRF_stage/reg_bank/n993 ,
         \iRF_stage/reg_bank/n992 , \iRF_stage/reg_bank/n991 ,
         \iRF_stage/reg_bank/n990 , \iRF_stage/reg_bank/n989 ,
         \iRF_stage/reg_bank/n988 , \iRF_stage/reg_bank/n987 ,
         \iRF_stage/reg_bank/n986 , \iRF_stage/reg_bank/n985 ,
         \iRF_stage/reg_bank/n984 , \iRF_stage/reg_bank/n983 ,
         \iRF_stage/reg_bank/n982 , \iRF_stage/reg_bank/n981 ,
         \iRF_stage/reg_bank/n980 , \iRF_stage/reg_bank/n979 ,
         \iRF_stage/reg_bank/n978 , \iRF_stage/reg_bank/n977 ,
         \iRF_stage/reg_bank/n976 , \iRF_stage/reg_bank/n975 ,
         \iRF_stage/reg_bank/n974 , \iRF_stage/reg_bank/n973 ,
         \iRF_stage/reg_bank/n972 , \iRF_stage/reg_bank/n971 ,
         \iRF_stage/reg_bank/n970 , \iRF_stage/reg_bank/n969 ,
         \iRF_stage/reg_bank/n968 , \iRF_stage/reg_bank/n967 ,
         \iRF_stage/reg_bank/n966 , \iRF_stage/reg_bank/n965 ,
         \iRF_stage/reg_bank/n964 , \iRF_stage/reg_bank/n963 ,
         \iRF_stage/reg_bank/n962 , \iRF_stage/reg_bank/n961 ,
         \iRF_stage/reg_bank/n960 , \iRF_stage/reg_bank/n959 ,
         \iRF_stage/reg_bank/n958 , \iRF_stage/reg_bank/n957 ,
         \iRF_stage/reg_bank/n956 , \iRF_stage/reg_bank/n955 ,
         \iRF_stage/reg_bank/n954 , \iRF_stage/reg_bank/n953 ,
         \iRF_stage/reg_bank/n952 , \iRF_stage/reg_bank/n951 ,
         \iRF_stage/reg_bank/n950 , \iRF_stage/reg_bank/n949 ,
         \iRF_stage/reg_bank/n948 , \iRF_stage/reg_bank/n947 ,
         \iRF_stage/reg_bank/n946 , \iRF_stage/reg_bank/n945 ,
         \iRF_stage/reg_bank/n944 , \iRF_stage/reg_bank/n943 ,
         \iRF_stage/reg_bank/n942 , \iRF_stage/reg_bank/n941 ,
         \iRF_stage/reg_bank/n940 , \iRF_stage/reg_bank/n939 ,
         \iRF_stage/reg_bank/n938 , \iRF_stage/reg_bank/n937 ,
         \iRF_stage/reg_bank/n936 , \iRF_stage/reg_bank/n935 ,
         \iRF_stage/reg_bank/n934 , \iRF_stage/reg_bank/n933 ,
         \iRF_stage/reg_bank/n932 , \iRF_stage/reg_bank/n931 ,
         \iRF_stage/reg_bank/n930 , \iRF_stage/reg_bank/n929 ,
         \iRF_stage/reg_bank/n928 , \iRF_stage/reg_bank/n927 ,
         \iRF_stage/reg_bank/n926 , \iRF_stage/reg_bank/n925 ,
         \iRF_stage/reg_bank/n924 , \iRF_stage/reg_bank/n923 ,
         \iRF_stage/reg_bank/n922 , \iRF_stage/reg_bank/n921 ,
         \iRF_stage/reg_bank/n920 , \iRF_stage/reg_bank/n919 ,
         \iRF_stage/reg_bank/n918 , \iRF_stage/reg_bank/n917 ,
         \iRF_stage/reg_bank/n916 , \iRF_stage/reg_bank/n915 ,
         \iRF_stage/reg_bank/n914 , \iRF_stage/reg_bank/n913 ,
         \iRF_stage/reg_bank/n912 , \iRF_stage/reg_bank/n911 ,
         \iRF_stage/reg_bank/n910 , \iRF_stage/reg_bank/n909 ,
         \iRF_stage/reg_bank/n908 , \iRF_stage/reg_bank/n907 ,
         \iRF_stage/reg_bank/n906 , \iRF_stage/reg_bank/n905 ,
         \iRF_stage/reg_bank/n904 , \iRF_stage/reg_bank/n903 ,
         \iRF_stage/reg_bank/n902 , \iRF_stage/reg_bank/n901 ,
         \iRF_stage/reg_bank/n900 , \iRF_stage/reg_bank/n899 ,
         \iRF_stage/reg_bank/n898 , \iRF_stage/reg_bank/n897 ,
         \iRF_stage/reg_bank/n896 , \iRF_stage/reg_bank/n895 ,
         \iRF_stage/reg_bank/n894 , \iRF_stage/reg_bank/n893 ,
         \iRF_stage/reg_bank/n892 , \iRF_stage/reg_bank/n891 ,
         \iRF_stage/reg_bank/n890 , \iRF_stage/reg_bank/n889 ,
         \iRF_stage/reg_bank/n888 , \iRF_stage/reg_bank/n887 ,
         \iRF_stage/reg_bank/n886 , \iRF_stage/reg_bank/n885 ,
         \iRF_stage/reg_bank/n884 , \iRF_stage/reg_bank/n883 ,
         \iRF_stage/reg_bank/n882 , \iRF_stage/reg_bank/n881 ,
         \iRF_stage/reg_bank/n880 , \iRF_stage/reg_bank/n879 ,
         \iRF_stage/reg_bank/n878 , \iRF_stage/reg_bank/n877 ,
         \iRF_stage/reg_bank/n876 , \iRF_stage/reg_bank/n875 ,
         \iRF_stage/reg_bank/n874 , \iRF_stage/reg_bank/n873 ,
         \iRF_stage/reg_bank/n872 , \iRF_stage/reg_bank/n871 ,
         \iRF_stage/reg_bank/n870 , \iRF_stage/reg_bank/n869 ,
         \iRF_stage/reg_bank/n868 , \iRF_stage/reg_bank/n867 ,
         \iRF_stage/reg_bank/n866 , \iRF_stage/reg_bank/n865 ,
         \iRF_stage/reg_bank/n864 , \iRF_stage/reg_bank/n863 ,
         \iRF_stage/reg_bank/n862 , \iRF_stage/reg_bank/n861 ,
         \iRF_stage/reg_bank/n860 , \iRF_stage/reg_bank/n859 ,
         \iRF_stage/reg_bank/n858 , \iRF_stage/reg_bank/n857 ,
         \iRF_stage/reg_bank/n856 , \iRF_stage/reg_bank/n855 ,
         \iRF_stage/reg_bank/n854 , \iRF_stage/reg_bank/n853 ,
         \iRF_stage/reg_bank/n852 , \iRF_stage/reg_bank/n851 ,
         \iRF_stage/reg_bank/n850 , \iRF_stage/reg_bank/n849 ,
         \iRF_stage/reg_bank/n848 , \iRF_stage/reg_bank/n847 ,
         \iRF_stage/reg_bank/n846 , \iRF_stage/reg_bank/n845 ,
         \iRF_stage/reg_bank/n844 , \iRF_stage/reg_bank/n843 ,
         \iRF_stage/reg_bank/n842 , \iRF_stage/reg_bank/n841 ,
         \iRF_stage/reg_bank/n840 , \iRF_stage/reg_bank/n839 ,
         \iRF_stage/reg_bank/n838 , \iRF_stage/reg_bank/n837 ,
         \iRF_stage/reg_bank/n836 , \iRF_stage/reg_bank/n835 ,
         \iRF_stage/reg_bank/n834 , \iRF_stage/reg_bank/n833 ,
         \iRF_stage/reg_bank/n832 , \iRF_stage/reg_bank/n831 ,
         \iRF_stage/reg_bank/n830 , \iRF_stage/reg_bank/n829 ,
         \iRF_stage/reg_bank/n828 , \iRF_stage/reg_bank/n827 ,
         \iRF_stage/reg_bank/n826 , \iRF_stage/reg_bank/n825 ,
         \iRF_stage/reg_bank/n824 , \iRF_stage/reg_bank/n823 ,
         \iRF_stage/reg_bank/n822 , \iRF_stage/reg_bank/n821 ,
         \iRF_stage/reg_bank/n820 , \iRF_stage/reg_bank/n819 ,
         \iRF_stage/reg_bank/n818 , \iRF_stage/reg_bank/n817 ,
         \iRF_stage/reg_bank/n816 , \iRF_stage/reg_bank/n815 ,
         \iRF_stage/reg_bank/n814 , \iRF_stage/reg_bank/n813 ,
         \iRF_stage/reg_bank/n812 , \iRF_stage/reg_bank/n811 ,
         \iRF_stage/reg_bank/n810 , \iRF_stage/reg_bank/n809 ,
         \iRF_stage/reg_bank/n808 , \iRF_stage/reg_bank/n807 ,
         \iRF_stage/reg_bank/n806 , \iRF_stage/reg_bank/n805 ,
         \iRF_stage/reg_bank/n804 , \iRF_stage/reg_bank/n803 ,
         \iRF_stage/reg_bank/n802 , \iRF_stage/reg_bank/n801 ,
         \iRF_stage/reg_bank/n800 , \iRF_stage/reg_bank/n799 ,
         \iRF_stage/reg_bank/n798 , \iRF_stage/reg_bank/n797 ,
         \iRF_stage/reg_bank/n796 , \iRF_stage/reg_bank/n795 ,
         \iRF_stage/reg_bank/n794 , \iRF_stage/reg_bank/n793 ,
         \iRF_stage/reg_bank/n792 , \iRF_stage/reg_bank/n791 ,
         \iRF_stage/reg_bank/n790 , \iRF_stage/reg_bank/n789 ,
         \iRF_stage/reg_bank/n788 , \iRF_stage/reg_bank/n787 ,
         \iRF_stage/reg_bank/n786 , \iRF_stage/reg_bank/n785 ,
         \iRF_stage/reg_bank/n784 , \iRF_stage/reg_bank/n783 ,
         \iRF_stage/reg_bank/n782 , \iRF_stage/reg_bank/n781 ,
         \iRF_stage/reg_bank/n780 , \iRF_stage/reg_bank/n779 ,
         \iRF_stage/reg_bank/n778 , \iRF_stage/reg_bank/n777 ,
         \iRF_stage/reg_bank/n776 , \iRF_stage/reg_bank/n775 ,
         \iRF_stage/reg_bank/n774 , \iRF_stage/reg_bank/n773 ,
         \iRF_stage/reg_bank/n772 , \iRF_stage/reg_bank/n771 ,
         \iRF_stage/reg_bank/n770 , \iRF_stage/reg_bank/n769 ,
         \iRF_stage/reg_bank/n768 , \iRF_stage/reg_bank/n767 ,
         \iRF_stage/reg_bank/n766 , \iRF_stage/reg_bank/n765 ,
         \iRF_stage/reg_bank/n764 , \iRF_stage/reg_bank/n763 ,
         \iRF_stage/reg_bank/n762 , \iRF_stage/reg_bank/n761 ,
         \iRF_stage/reg_bank/n760 , \iRF_stage/reg_bank/n759 ,
         \iRF_stage/reg_bank/n758 , \iRF_stage/reg_bank/n757 ,
         \iRF_stage/reg_bank/n756 , \iRF_stage/reg_bank/n755 ,
         \iRF_stage/reg_bank/n754 , \iRF_stage/reg_bank/n753 ,
         \iRF_stage/reg_bank/n752 , \iRF_stage/reg_bank/n751 ,
         \iRF_stage/reg_bank/n750 , \iRF_stage/reg_bank/n749 ,
         \iRF_stage/reg_bank/n748 , \iRF_stage/reg_bank/n747 ,
         \iRF_stage/reg_bank/n746 , \iRF_stage/reg_bank/n745 ,
         \iRF_stage/reg_bank/n744 , \iRF_stage/reg_bank/n743 ,
         \iRF_stage/reg_bank/n742 , \iRF_stage/reg_bank/n741 ,
         \iRF_stage/reg_bank/n740 , \iRF_stage/reg_bank/n739 ,
         \iRF_stage/reg_bank/n738 , \iRF_stage/reg_bank/n737 ,
         \iRF_stage/reg_bank/n736 , \iRF_stage/reg_bank/n735 ,
         \iRF_stage/reg_bank/n734 , \iRF_stage/reg_bank/n733 ,
         \iRF_stage/reg_bank/n732 , \iRF_stage/reg_bank/n731 ,
         \iRF_stage/reg_bank/n730 , \iRF_stage/reg_bank/n729 ,
         \iRF_stage/reg_bank/n728 , \iRF_stage/reg_bank/n727 ,
         \iRF_stage/reg_bank/n726 , \iRF_stage/reg_bank/n725 ,
         \iRF_stage/reg_bank/n724 , \iRF_stage/reg_bank/n723 ,
         \iRF_stage/reg_bank/n722 , \iRF_stage/reg_bank/n721 ,
         \iRF_stage/reg_bank/n720 , \iRF_stage/reg_bank/n719 ,
         \iRF_stage/reg_bank/n718 , \iRF_stage/reg_bank/n717 ,
         \iRF_stage/reg_bank/n716 , \iRF_stage/reg_bank/n715 ,
         \iRF_stage/reg_bank/n714 , \iRF_stage/reg_bank/n713 ,
         \iRF_stage/reg_bank/n712 , \iRF_stage/reg_bank/n711 ,
         \iRF_stage/reg_bank/n710 , \iRF_stage/reg_bank/n709 ,
         \iRF_stage/reg_bank/n708 , \iRF_stage/reg_bank/n707 ,
         \iRF_stage/reg_bank/n706 , \iRF_stage/reg_bank/n705 ,
         \iRF_stage/reg_bank/n704 , \iRF_stage/reg_bank/n703 ,
         \iRF_stage/reg_bank/n702 , \iRF_stage/reg_bank/n701 ,
         \iRF_stage/reg_bank/n700 , \iRF_stage/reg_bank/n699 ,
         \iRF_stage/reg_bank/n698 , \iRF_stage/reg_bank/n697 ,
         \iRF_stage/reg_bank/n696 , \iRF_stage/reg_bank/n695 ,
         \iRF_stage/reg_bank/n694 , \iRF_stage/reg_bank/n693 ,
         \iRF_stage/reg_bank/n692 , \iRF_stage/reg_bank/n691 ,
         \iRF_stage/reg_bank/n690 , \iRF_stage/reg_bank/n689 ,
         \iRF_stage/reg_bank/n688 , \iRF_stage/reg_bank/n687 ,
         \iRF_stage/reg_bank/n686 , \iRF_stage/reg_bank/n685 ,
         \iRF_stage/reg_bank/n684 , \iRF_stage/reg_bank/n683 ,
         \iRF_stage/reg_bank/n682 , \iRF_stage/reg_bank/n681 ,
         \iRF_stage/reg_bank/n680 , \iRF_stage/reg_bank/n679 ,
         \iRF_stage/reg_bank/n678 , \iRF_stage/reg_bank/n677 ,
         \iRF_stage/reg_bank/n676 , \iRF_stage/reg_bank/n675 ,
         \iRF_stage/reg_bank/n674 , \iRF_stage/reg_bank/n673 ,
         \iRF_stage/reg_bank/n672 , \iRF_stage/reg_bank/n671 ,
         \iRF_stage/reg_bank/n670 , \iRF_stage/reg_bank/n669 ,
         \iRF_stage/reg_bank/n668 , \iRF_stage/reg_bank/n667 ,
         \iRF_stage/reg_bank/n666 , \iRF_stage/reg_bank/n665 ,
         \iRF_stage/reg_bank/n664 , \iRF_stage/reg_bank/n663 ,
         \iRF_stage/reg_bank/n662 , \iRF_stage/reg_bank/n661 ,
         \iRF_stage/reg_bank/n660 , \iRF_stage/reg_bank/n659 ,
         \iRF_stage/reg_bank/n658 , \iRF_stage/reg_bank/n657 ,
         \iRF_stage/reg_bank/n656 , \iRF_stage/reg_bank/n655 ,
         \iRF_stage/reg_bank/n654 , \iRF_stage/reg_bank/n653 ,
         \iRF_stage/reg_bank/n652 , \iRF_stage/reg_bank/n651 ,
         \iRF_stage/reg_bank/n650 , \iRF_stage/reg_bank/n649 ,
         \iRF_stage/reg_bank/n648 , \iRF_stage/reg_bank/n647 ,
         \iRF_stage/reg_bank/n646 , \iRF_stage/reg_bank/n645 ,
         \iRF_stage/reg_bank/n644 , \iRF_stage/reg_bank/n643 ,
         \iRF_stage/reg_bank/n642 , \iRF_stage/reg_bank/n641 ,
         \iRF_stage/reg_bank/n640 , \iRF_stage/reg_bank/n639 ,
         \iRF_stage/reg_bank/n638 , \iRF_stage/reg_bank/n637 ,
         \iRF_stage/reg_bank/n636 , \iRF_stage/reg_bank/n635 ,
         \iRF_stage/reg_bank/n634 , \iRF_stage/reg_bank/n633 ,
         \iRF_stage/reg_bank/n632 , \iRF_stage/reg_bank/n631 ,
         \iRF_stage/reg_bank/n630 , \iRF_stage/reg_bank/n629 ,
         \iRF_stage/reg_bank/n628 , \iRF_stage/reg_bank/n627 ,
         \iRF_stage/reg_bank/n626 , \iRF_stage/reg_bank/n625 ,
         \iRF_stage/reg_bank/n624 , \iRF_stage/reg_bank/n623 ,
         \iRF_stage/reg_bank/n622 , \iRF_stage/reg_bank/n621 ,
         \iRF_stage/reg_bank/n620 , \iRF_stage/reg_bank/n619 ,
         \iRF_stage/reg_bank/n618 , \iRF_stage/reg_bank/n617 ,
         \iRF_stage/reg_bank/n616 , \iRF_stage/reg_bank/n615 ,
         \iRF_stage/reg_bank/n614 , \iRF_stage/reg_bank/n613 ,
         \iRF_stage/reg_bank/n612 , \iRF_stage/reg_bank/n611 ,
         \iRF_stage/reg_bank/n610 , \iRF_stage/reg_bank/n609 ,
         \iRF_stage/reg_bank/n608 , \iRF_stage/reg_bank/n607 ,
         \iRF_stage/reg_bank/n606 , \iRF_stage/reg_bank/n605 ,
         \iRF_stage/reg_bank/n604 , \iRF_stage/reg_bank/n603 ,
         \iRF_stage/reg_bank/n602 , \iRF_stage/reg_bank/n601 ,
         \iRF_stage/reg_bank/n600 , \iRF_stage/reg_bank/n599 ,
         \iRF_stage/reg_bank/n598 , \iRF_stage/reg_bank/n597 ,
         \iRF_stage/reg_bank/n596 , \iRF_stage/reg_bank/n595 ,
         \iRF_stage/reg_bank/n594 , \iRF_stage/reg_bank/n593 ,
         \iRF_stage/reg_bank/n592 , \iRF_stage/reg_bank/n591 ,
         \iRF_stage/reg_bank/n590 , \iRF_stage/reg_bank/n589 ,
         \iRF_stage/reg_bank/n588 , \iRF_stage/reg_bank/n587 ,
         \iRF_stage/reg_bank/n586 , \iRF_stage/reg_bank/n585 ,
         \iRF_stage/reg_bank/n584 , \iRF_stage/reg_bank/n583 ,
         \iRF_stage/reg_bank/n582 , \iRF_stage/reg_bank/n581 ,
         \iRF_stage/reg_bank/n580 , \iRF_stage/reg_bank/n579 ,
         \iRF_stage/reg_bank/n578 , \iRF_stage/reg_bank/n577 ,
         \iRF_stage/reg_bank/n576 , \iRF_stage/reg_bank/n575 ,
         \iRF_stage/reg_bank/n574 , \iRF_stage/reg_bank/n573 ,
         \iRF_stage/reg_bank/n572 , \iRF_stage/reg_bank/n571 ,
         \iRF_stage/reg_bank/n570 , \iRF_stage/reg_bank/n569 ,
         \iRF_stage/reg_bank/n568 , \iRF_stage/reg_bank/n567 ,
         \iRF_stage/reg_bank/n566 , \iRF_stage/reg_bank/n565 ,
         \iRF_stage/reg_bank/n564 , \iRF_stage/reg_bank/n563 ,
         \iRF_stage/reg_bank/n562 , \iRF_stage/reg_bank/n561 ,
         \iRF_stage/reg_bank/n560 , \iRF_stage/reg_bank/n559 ,
         \iRF_stage/reg_bank/n558 , \iRF_stage/reg_bank/n557 ,
         \iRF_stage/reg_bank/n556 , \iRF_stage/reg_bank/n555 ,
         \iRF_stage/reg_bank/n554 , \iRF_stage/reg_bank/n553 ,
         \iRF_stage/reg_bank/n552 , \iRF_stage/reg_bank/n551 ,
         \iRF_stage/reg_bank/n550 , \iRF_stage/reg_bank/n549 ,
         \iRF_stage/reg_bank/n548 , \iRF_stage/reg_bank/n547 ,
         \iRF_stage/reg_bank/n546 , \iRF_stage/reg_bank/n545 ,
         \iRF_stage/reg_bank/n544 , \iRF_stage/reg_bank/n543 ,
         \iRF_stage/reg_bank/n542 , \iRF_stage/reg_bank/n541 ,
         \iRF_stage/reg_bank/n540 , \iRF_stage/reg_bank/n539 ,
         \iRF_stage/reg_bank/n538 , \iRF_stage/reg_bank/n537 ,
         \iRF_stage/reg_bank/n536 , \iRF_stage/reg_bank/n535 ,
         \iRF_stage/reg_bank/n534 , \iRF_stage/reg_bank/n533 ,
         \iRF_stage/reg_bank/n532 , \iRF_stage/reg_bank/n531 ,
         \iRF_stage/reg_bank/n530 , \iRF_stage/reg_bank/n529 ,
         \iRF_stage/reg_bank/n528 , \iRF_stage/reg_bank/n527 ,
         \iRF_stage/reg_bank/n526 , \iRF_stage/reg_bank/n525 ,
         \iRF_stage/reg_bank/n524 , \iRF_stage/reg_bank/n523 ,
         \iRF_stage/reg_bank/n522 , \iRF_stage/reg_bank/n521 ,
         \iRF_stage/reg_bank/n520 , \iRF_stage/reg_bank/n519 ,
         \iRF_stage/reg_bank/n518 , \iRF_stage/reg_bank/n517 ,
         \iRF_stage/reg_bank/n516 , \iRF_stage/reg_bank/n515 ,
         \iRF_stage/reg_bank/n514 , \iRF_stage/reg_bank/n513 ,
         \iRF_stage/reg_bank/n512 , \iRF_stage/reg_bank/n511 ,
         \iRF_stage/reg_bank/n510 , \iRF_stage/reg_bank/n509 ,
         \iRF_stage/reg_bank/n508 , \iRF_stage/reg_bank/n507 ,
         \iRF_stage/reg_bank/n506 , \iRF_stage/reg_bank/n505 ,
         \iRF_stage/reg_bank/n504 , \iRF_stage/reg_bank/n503 ,
         \iRF_stage/reg_bank/n502 , \iRF_stage/reg_bank/n501 ,
         \iRF_stage/reg_bank/n500 , \iRF_stage/reg_bank/n499 ,
         \iRF_stage/reg_bank/n498 , \iRF_stage/reg_bank/n497 ,
         \iRF_stage/reg_bank/n496 , \iRF_stage/reg_bank/n495 ,
         \iRF_stage/reg_bank/n494 , \iRF_stage/reg_bank/n493 ,
         \iRF_stage/reg_bank/n492 , \iRF_stage/reg_bank/n491 ,
         \iRF_stage/reg_bank/n490 , \iRF_stage/reg_bank/n489 ,
         \iRF_stage/reg_bank/n488 , \iRF_stage/reg_bank/n487 ,
         \iRF_stage/reg_bank/n486 , \iRF_stage/reg_bank/n485 ,
         \iRF_stage/reg_bank/n484 , \iRF_stage/reg_bank/n483 ,
         \iRF_stage/reg_bank/n482 , \iRF_stage/reg_bank/n481 ,
         \iRF_stage/reg_bank/n480 , \iRF_stage/reg_bank/n479 ,
         \iRF_stage/reg_bank/n478 , \iRF_stage/reg_bank/n477 ,
         \iRF_stage/reg_bank/n476 , \iRF_stage/reg_bank/n475 ,
         \iRF_stage/reg_bank/n474 , \iRF_stage/reg_bank/n473 ,
         \iRF_stage/reg_bank/n472 , \iRF_stage/reg_bank/n471 ,
         \iRF_stage/reg_bank/n470 , \iRF_stage/reg_bank/n469 ,
         \iRF_stage/reg_bank/n468 , \iRF_stage/reg_bank/n467 ,
         \iRF_stage/reg_bank/n466 , \iRF_stage/reg_bank/n465 ,
         \iRF_stage/reg_bank/n464 , \iRF_stage/reg_bank/n463 ,
         \iRF_stage/reg_bank/n462 , \iRF_stage/reg_bank/n461 ,
         \iRF_stage/reg_bank/n460 , \iRF_stage/reg_bank/n459 ,
         \iRF_stage/reg_bank/n458 , \iRF_stage/reg_bank/n457 ,
         \iRF_stage/reg_bank/n456 , \iRF_stage/reg_bank/n455 ,
         \iRF_stage/reg_bank/n454 , \iRF_stage/reg_bank/n453 ,
         \iRF_stage/reg_bank/n452 , \iRF_stage/reg_bank/n451 ,
         \iRF_stage/reg_bank/n450 , \iRF_stage/reg_bank/n449 ,
         \iRF_stage/reg_bank/n448 , \iRF_stage/reg_bank/n447 ,
         \iRF_stage/reg_bank/n446 , \iRF_stage/reg_bank/n445 ,
         \iRF_stage/reg_bank/n444 , \iRF_stage/reg_bank/n443 ,
         \iRF_stage/reg_bank/n442 , \iRF_stage/reg_bank/n441 ,
         \iRF_stage/reg_bank/n440 , \iRF_stage/reg_bank/n439 ,
         \iRF_stage/reg_bank/n438 , \iRF_stage/reg_bank/n437 ,
         \iRF_stage/reg_bank/n436 , \iRF_stage/reg_bank/n435 ,
         \iRF_stage/reg_bank/n434 , \iRF_stage/reg_bank/n433 ,
         \iRF_stage/reg_bank/n432 , \iRF_stage/reg_bank/n431 ,
         \iRF_stage/reg_bank/n430 , \iRF_stage/reg_bank/n429 ,
         \iRF_stage/reg_bank/n428 , \iRF_stage/reg_bank/n427 ,
         \iRF_stage/reg_bank/n426 , \iRF_stage/reg_bank/n425 ,
         \iRF_stage/reg_bank/n424 , \iRF_stage/reg_bank/n423 ,
         \iRF_stage/reg_bank/n422 , \iRF_stage/reg_bank/n421 ,
         \iRF_stage/reg_bank/n420 , \iRF_stage/reg_bank/n419 ,
         \iRF_stage/reg_bank/n418 , \iRF_stage/reg_bank/n417 ,
         \iRF_stage/reg_bank/n416 , \iRF_stage/reg_bank/n415 ,
         \iRF_stage/reg_bank/n414 , \iRF_stage/reg_bank/n413 ,
         \iRF_stage/reg_bank/n412 , \iRF_stage/reg_bank/n411 ,
         \iRF_stage/reg_bank/n410 , \iRF_stage/reg_bank/n409 ,
         \iRF_stage/reg_bank/n408 , \iRF_stage/reg_bank/n407 ,
         \iRF_stage/reg_bank/n406 , \iRF_stage/reg_bank/n405 ,
         \iRF_stage/reg_bank/n404 , \iRF_stage/reg_bank/n403 ,
         \iRF_stage/reg_bank/n402 , \iRF_stage/reg_bank/n401 ,
         \iRF_stage/reg_bank/n400 , \iRF_stage/reg_bank/n399 ,
         \iRF_stage/reg_bank/n398 , \iRF_stage/reg_bank/n397 ,
         \iRF_stage/reg_bank/n396 , \iRF_stage/reg_bank/n395 ,
         \iRF_stage/reg_bank/n394 , \iRF_stage/reg_bank/n393 ,
         \iRF_stage/reg_bank/n392 , \iRF_stage/reg_bank/n391 ,
         \iRF_stage/reg_bank/n390 , \iRF_stage/reg_bank/n389 ,
         \iRF_stage/reg_bank/n388 , \iRF_stage/reg_bank/n387 ,
         \iRF_stage/reg_bank/n386 , \iRF_stage/reg_bank/n385 ,
         \iRF_stage/reg_bank/n384 , \iRF_stage/reg_bank/n383 ,
         \iRF_stage/reg_bank/n382 , \iRF_stage/reg_bank/n381 ,
         \iRF_stage/reg_bank/n380 , \iRF_stage/reg_bank/n379 ,
         \iRF_stage/reg_bank/n378 , \iRF_stage/reg_bank/n377 ,
         \iRF_stage/reg_bank/n376 , \iRF_stage/reg_bank/n375 ,
         \iRF_stage/reg_bank/n374 , \iRF_stage/reg_bank/n373 ,
         \iRF_stage/reg_bank/n372 , \iRF_stage/reg_bank/n371 ,
         \iRF_stage/reg_bank/n370 , \iRF_stage/reg_bank/n369 ,
         \iRF_stage/reg_bank/n368 , \iRF_stage/reg_bank/n367 ,
         \iRF_stage/reg_bank/n366 , \iRF_stage/reg_bank/n365 ,
         \iRF_stage/reg_bank/n364 , \iRF_stage/reg_bank/n363 ,
         \iRF_stage/reg_bank/n362 , \iRF_stage/reg_bank/n361 ,
         \iRF_stage/reg_bank/n360 , \iRF_stage/reg_bank/n359 ,
         \iRF_stage/reg_bank/n358 , \iRF_stage/reg_bank/n357 ,
         \iRF_stage/reg_bank/n356 , \iRF_stage/reg_bank/n355 ,
         \iRF_stage/reg_bank/n354 , \iRF_stage/reg_bank/n353 ,
         \iRF_stage/reg_bank/n352 , \iRF_stage/reg_bank/n351 ,
         \iRF_stage/reg_bank/n350 , \iRF_stage/reg_bank/n349 ,
         \iRF_stage/reg_bank/n348 , \iRF_stage/reg_bank/n347 ,
         \iRF_stage/reg_bank/n346 , \iRF_stage/reg_bank/n345 ,
         \iRF_stage/reg_bank/n344 , \iRF_stage/reg_bank/n343 ,
         \iRF_stage/reg_bank/n342 , \iRF_stage/reg_bank/n341 ,
         \iRF_stage/reg_bank/n340 , \iRF_stage/reg_bank/n339 ,
         \iRF_stage/reg_bank/n338 , \iRF_stage/reg_bank/n337 ,
         \iRF_stage/reg_bank/n336 , \iRF_stage/reg_bank/n335 ,
         \iRF_stage/reg_bank/n334 , \iRF_stage/reg_bank/n333 ,
         \iRF_stage/reg_bank/n332 , \iRF_stage/reg_bank/n331 ,
         \iRF_stage/reg_bank/n330 , \iRF_stage/reg_bank/n329 ,
         \iRF_stage/reg_bank/n328 , \iRF_stage/reg_bank/n327 ,
         \iRF_stage/reg_bank/n326 , \iRF_stage/reg_bank/n325 ,
         \iRF_stage/reg_bank/n324 , \iRF_stage/reg_bank/n323 ,
         \iRF_stage/reg_bank/n322 , \iRF_stage/reg_bank/n321 ,
         \iRF_stage/reg_bank/n320 , \iRF_stage/reg_bank/n319 ,
         \iRF_stage/reg_bank/n318 , \iRF_stage/reg_bank/n317 ,
         \iRF_stage/reg_bank/n316 , \iRF_stage/reg_bank/n315 ,
         \iRF_stage/reg_bank/n314 , \iRF_stage/reg_bank/n313 ,
         \iRF_stage/reg_bank/n312 , \iRF_stage/reg_bank/n311 ,
         \iRF_stage/reg_bank/n310 , \iRF_stage/reg_bank/n309 ,
         \iRF_stage/reg_bank/n308 , \iRF_stage/reg_bank/n307 ,
         \iRF_stage/reg_bank/n306 , \iRF_stage/reg_bank/n305 ,
         \iRF_stage/reg_bank/n304 , \iRF_stage/reg_bank/n303 ,
         \iRF_stage/reg_bank/n302 , \iRF_stage/reg_bank/n301 ,
         \iRF_stage/reg_bank/n300 , \iRF_stage/reg_bank/n299 ,
         \iRF_stage/reg_bank/n298 , \iRF_stage/reg_bank/n297 ,
         \iRF_stage/reg_bank/n296 , \iRF_stage/reg_bank/n295 ,
         \iRF_stage/reg_bank/n294 , \iRF_stage/reg_bank/n293 ,
         \iRF_stage/reg_bank/n292 , \iRF_stage/reg_bank/n291 ,
         \iRF_stage/reg_bank/n290 , \iRF_stage/reg_bank/n289 ,
         \iRF_stage/reg_bank/n288 , \iRF_stage/reg_bank/n287 ,
         \iRF_stage/reg_bank/n286 , \iRF_stage/reg_bank/n285 ,
         \iRF_stage/reg_bank/n284 , \iRF_stage/reg_bank/n283 ,
         \iRF_stage/reg_bank/n282 , \iRF_stage/reg_bank/n281 ,
         \iRF_stage/reg_bank/n280 , \iRF_stage/reg_bank/n279 ,
         \iRF_stage/reg_bank/n278 , \iRF_stage/reg_bank/n277 ,
         \iRF_stage/reg_bank/n276 , \iRF_stage/reg_bank/n275 ,
         \iRF_stage/reg_bank/n274 , \iRF_stage/reg_bank/n273 ,
         \iRF_stage/reg_bank/n272 , \iRF_stage/reg_bank/n271 ,
         \iRF_stage/reg_bank/n270 , \iRF_stage/reg_bank/n269 ,
         \iRF_stage/reg_bank/n268 , \iRF_stage/reg_bank/n267 ,
         \iRF_stage/reg_bank/n266 , \iRF_stage/reg_bank/n265 ,
         \iRF_stage/reg_bank/n264 , \iRF_stage/reg_bank/n263 ,
         \iRF_stage/reg_bank/n262 , \iRF_stage/reg_bank/n261 ,
         \iRF_stage/reg_bank/n260 , \iRF_stage/reg_bank/n259 ,
         \iRF_stage/reg_bank/n258 , \iRF_stage/reg_bank/n257 ,
         \iRF_stage/reg_bank/n256 , \iRF_stage/reg_bank/n255 ,
         \iRF_stage/reg_bank/n254 , \iRF_stage/reg_bank/n253 ,
         \iRF_stage/reg_bank/n252 , \iRF_stage/reg_bank/n251 ,
         \iRF_stage/reg_bank/n250 , \iRF_stage/reg_bank/n249 ,
         \iRF_stage/reg_bank/n248 , \iRF_stage/reg_bank/n247 ,
         \iRF_stage/reg_bank/n246 , \iRF_stage/reg_bank/n245 ,
         \iRF_stage/reg_bank/n244 , \iRF_stage/reg_bank/n243 ,
         \iRF_stage/reg_bank/n242 , \iRF_stage/reg_bank/n241 ,
         \iRF_stage/reg_bank/n240 , \iRF_stage/reg_bank/n239 ,
         \iRF_stage/reg_bank/n238 , \iRF_stage/reg_bank/n237 ,
         \iRF_stage/reg_bank/n236 , \iRF_stage/reg_bank/n235 ,
         \iRF_stage/reg_bank/n234 , \iRF_stage/reg_bank/n233 ,
         \iRF_stage/reg_bank/n232 , \iRF_stage/reg_bank/n231 ,
         \iRF_stage/reg_bank/n230 , \iRF_stage/reg_bank/n229 ,
         \iRF_stage/reg_bank/n228 , \iRF_stage/reg_bank/n227 ,
         \iRF_stage/reg_bank/n226 , \iRF_stage/reg_bank/n225 ,
         \iRF_stage/reg_bank/n224 , \iRF_stage/reg_bank/n223 ,
         \iRF_stage/reg_bank/n222 , \iRF_stage/reg_bank/n221 ,
         \iRF_stage/reg_bank/n220 , \iRF_stage/reg_bank/n219 ,
         \iRF_stage/reg_bank/n218 , \iRF_stage/reg_bank/n217 ,
         \iRF_stage/reg_bank/n216 , \iRF_stage/reg_bank/n215 ,
         \iRF_stage/reg_bank/n214 , \iRF_stage/reg_bank/n213 ,
         \iRF_stage/reg_bank/n212 , \iRF_stage/reg_bank/n211 ,
         \iRF_stage/reg_bank/n210 , \iRF_stage/reg_bank/n209 ,
         \iRF_stage/reg_bank/n208 , \iRF_stage/reg_bank/n207 ,
         \iRF_stage/reg_bank/n206 , \iRF_stage/reg_bank/n205 ,
         \iRF_stage/reg_bank/n204 , \iRF_stage/reg_bank/n203 ,
         \iRF_stage/reg_bank/n202 , \iRF_stage/reg_bank/n201 ,
         \iRF_stage/reg_bank/n200 , \iRF_stage/reg_bank/n199 ,
         \iRF_stage/reg_bank/n198 , \iRF_stage/reg_bank/n197 ,
         \iRF_stage/reg_bank/n196 , \iRF_stage/reg_bank/n195 ,
         \iRF_stage/reg_bank/n194 , \iRF_stage/reg_bank/n193 ,
         \iRF_stage/reg_bank/n192 , \iRF_stage/reg_bank/n191 ,
         \iRF_stage/reg_bank/n190 , \iRF_stage/reg_bank/n189 ,
         \iRF_stage/reg_bank/n188 , \iRF_stage/reg_bank/n187 ,
         \iRF_stage/reg_bank/n186 , \iRF_stage/reg_bank/n185 ,
         \iRF_stage/reg_bank/n184 , \iRF_stage/reg_bank/n183 ,
         \iRF_stage/reg_bank/n182 , \iRF_stage/reg_bank/n181 ,
         \iRF_stage/reg_bank/n180 , \iRF_stage/reg_bank/n179 ,
         \iRF_stage/reg_bank/n178 , \iRF_stage/reg_bank/n177 ,
         \iRF_stage/reg_bank/n176 , \iRF_stage/reg_bank/n175 ,
         \iRF_stage/reg_bank/n174 , \iRF_stage/reg_bank/n173 ,
         \iRF_stage/reg_bank/n172 , \iRF_stage/reg_bank/n171 ,
         \iRF_stage/reg_bank/n170 , \iRF_stage/reg_bank/n169 ,
         \iRF_stage/reg_bank/n168 , \iRF_stage/reg_bank/n167 ,
         \iRF_stage/reg_bank/n166 , \iRF_stage/reg_bank/n165 ,
         \iRF_stage/reg_bank/n164 , \iRF_stage/reg_bank/n163 ,
         \iRF_stage/reg_bank/n162 , \iRF_stage/reg_bank/n161 ,
         \iRF_stage/reg_bank/n160 , \iRF_stage/reg_bank/n159 ,
         \iRF_stage/reg_bank/n158 , \iRF_stage/reg_bank/n157 ,
         \iRF_stage/reg_bank/n156 , \iRF_stage/reg_bank/n155 ,
         \iRF_stage/reg_bank/n154 , \iRF_stage/reg_bank/n153 ,
         \iRF_stage/reg_bank/n152 , \iRF_stage/reg_bank/n151 ,
         \iRF_stage/reg_bank/n150 , \iRF_stage/reg_bank/n149 ,
         \iRF_stage/reg_bank/n148 , \iRF_stage/reg_bank/n147 ,
         \iRF_stage/reg_bank/n146 , \iRF_stage/reg_bank/n145 ,
         \iRF_stage/reg_bank/n144 , \iRF_stage/reg_bank/n143 ,
         \iRF_stage/reg_bank/n142 , \iRF_stage/reg_bank/n141 ,
         \iRF_stage/reg_bank/n140 , \iRF_stage/reg_bank/n139 ,
         \iRF_stage/reg_bank/n138 , \iRF_stage/reg_bank/N1120 ,
         \iRF_stage/reg_bank/N1119 , \iRF_stage/reg_bank/N1118 ,
         \iRF_stage/reg_bank/N1117 , \iRF_stage/reg_bank/N1116 ,
         \iRF_stage/reg_bank/N1115 , \iRF_stage/reg_bank/N1114 ,
         \iRF_stage/reg_bank/N1113 , \iRF_stage/reg_bank/N1112 ,
         \iRF_stage/reg_bank/N1111 , \iRF_stage/reg_bank/N1110 ,
         \iRF_stage/reg_bank/N1109 , \iRF_stage/reg_bank/N1108 ,
         \iRF_stage/reg_bank/N1107 , \iRF_stage/reg_bank/N1106 ,
         \iRF_stage/reg_bank/N1105 , \iRF_stage/reg_bank/N1104 ,
         \iRF_stage/reg_bank/N1103 , \iRF_stage/reg_bank/N1102 ,
         \iRF_stage/reg_bank/N1101 , \iRF_stage/reg_bank/N1100 ,
         \iRF_stage/reg_bank/N1099 , \iRF_stage/reg_bank/N1098 ,
         \iRF_stage/reg_bank/N1097 , \iRF_stage/reg_bank/N1096 ,
         \iRF_stage/reg_bank/N1095 , \iRF_stage/reg_bank/N1094 ,
         \iRF_stage/reg_bank/N1093 , \iRF_stage/reg_bank/N1092 ,
         \iRF_stage/reg_bank/N1091 , \iRF_stage/reg_bank/N1090 ,
         \iRF_stage/reg_bank/N1089 , \iRF_stage/reg_bank/N1083 ,
         \iRF_stage/reg_bank/N1082 , \iRF_stage/reg_bank/N1081 ,
         \iRF_stage/reg_bank/N1080 , \iRF_stage/reg_bank/N1079 ,
         \iRF_stage/reg_bank/N1078 , \iRF_stage/reg_bank/N1077 ,
         \iRF_stage/reg_bank/N1076 , \iRF_stage/reg_bank/N1075 ,
         \iRF_stage/reg_bank/N1074 , \iRF_stage/reg_bank/N1073 ,
         \iRF_stage/reg_bank/N1072 , \iRF_stage/reg_bank/N1071 ,
         \iRF_stage/reg_bank/N1070 , \iRF_stage/reg_bank/N1069 ,
         \iRF_stage/reg_bank/N1068 , \iRF_stage/reg_bank/N1067 ,
         \iRF_stage/reg_bank/N1066 , \iRF_stage/reg_bank/N1065 ,
         \iRF_stage/reg_bank/N1064 , \iRF_stage/reg_bank/N1063 ,
         \iRF_stage/reg_bank/N1062 , \iRF_stage/reg_bank/N1061 ,
         \iRF_stage/reg_bank/N1060 , \iRF_stage/reg_bank/N1059 ,
         \iRF_stage/reg_bank/N1058 , \iRF_stage/reg_bank/N1057 ,
         \iRF_stage/reg_bank/N1056 , \iRF_stage/reg_bank/N1055 ,
         \iRF_stage/reg_bank/N1054 , \iRF_stage/reg_bank/N1053 ,
         \iRF_stage/reg_bank/N1052 , \iRF_stage/reg_bank/reg_bank[0] ,
         \iRF_stage/reg_bank/reg_bank[1] , \iRF_stage/reg_bank/reg_bank[2] ,
         \iRF_stage/reg_bank/reg_bank[3] , \iRF_stage/reg_bank/reg_bank[4] ,
         \iRF_stage/reg_bank/reg_bank[5] , \iRF_stage/reg_bank/reg_bank[6] ,
         \iRF_stage/reg_bank/reg_bank[7] , \iRF_stage/reg_bank/reg_bank[8] ,
         \iRF_stage/reg_bank/reg_bank[9] , \iRF_stage/reg_bank/reg_bank[10] ,
         \iRF_stage/reg_bank/reg_bank[11] , \iRF_stage/reg_bank/reg_bank[12] ,
         \iRF_stage/reg_bank/reg_bank[13] , \iRF_stage/reg_bank/reg_bank[14] ,
         \iRF_stage/reg_bank/reg_bank[15] , \iRF_stage/reg_bank/reg_bank[16] ,
         \iRF_stage/reg_bank/reg_bank[17] , \iRF_stage/reg_bank/reg_bank[18] ,
         \iRF_stage/reg_bank/reg_bank[19] , \iRF_stage/reg_bank/reg_bank[20] ,
         \iRF_stage/reg_bank/reg_bank[21] , \iRF_stage/reg_bank/reg_bank[22] ,
         \iRF_stage/reg_bank/reg_bank[23] , \iRF_stage/reg_bank/reg_bank[24] ,
         \iRF_stage/reg_bank/reg_bank[25] , \iRF_stage/reg_bank/reg_bank[26] ,
         \iRF_stage/reg_bank/reg_bank[27] , \iRF_stage/reg_bank/reg_bank[28] ,
         \iRF_stage/reg_bank/reg_bank[29] , \iRF_stage/reg_bank/reg_bank[30] ,
         \iRF_stage/reg_bank/reg_bank[31] , \iRF_stage/reg_bank/reg_bank[32] ,
         \iRF_stage/reg_bank/reg_bank[33] , \iRF_stage/reg_bank/reg_bank[34] ,
         \iRF_stage/reg_bank/reg_bank[35] , \iRF_stage/reg_bank/reg_bank[36] ,
         \iRF_stage/reg_bank/reg_bank[37] , \iRF_stage/reg_bank/reg_bank[38] ,
         \iRF_stage/reg_bank/reg_bank[39] , \iRF_stage/reg_bank/reg_bank[40] ,
         \iRF_stage/reg_bank/reg_bank[41] , \iRF_stage/reg_bank/reg_bank[42] ,
         \iRF_stage/reg_bank/reg_bank[43] , \iRF_stage/reg_bank/reg_bank[44] ,
         \iRF_stage/reg_bank/reg_bank[45] , \iRF_stage/reg_bank/reg_bank[46] ,
         \iRF_stage/reg_bank/reg_bank[47] , \iRF_stage/reg_bank/reg_bank[48] ,
         \iRF_stage/reg_bank/reg_bank[49] , \iRF_stage/reg_bank/reg_bank[50] ,
         \iRF_stage/reg_bank/reg_bank[51] , \iRF_stage/reg_bank/reg_bank[52] ,
         \iRF_stage/reg_bank/reg_bank[53] , \iRF_stage/reg_bank/reg_bank[54] ,
         \iRF_stage/reg_bank/reg_bank[55] , \iRF_stage/reg_bank/reg_bank[56] ,
         \iRF_stage/reg_bank/reg_bank[57] , \iRF_stage/reg_bank/reg_bank[58] ,
         \iRF_stage/reg_bank/reg_bank[59] , \iRF_stage/reg_bank/reg_bank[60] ,
         \iRF_stage/reg_bank/reg_bank[61] , \iRF_stage/reg_bank/reg_bank[62] ,
         \iRF_stage/reg_bank/reg_bank[63] , \iRF_stage/reg_bank/reg_bank[64] ,
         \iRF_stage/reg_bank/reg_bank[65] , \iRF_stage/reg_bank/reg_bank[66] ,
         \iRF_stage/reg_bank/reg_bank[67] , \iRF_stage/reg_bank/reg_bank[68] ,
         \iRF_stage/reg_bank/reg_bank[69] , \iRF_stage/reg_bank/reg_bank[70] ,
         \iRF_stage/reg_bank/reg_bank[71] , \iRF_stage/reg_bank/reg_bank[72] ,
         \iRF_stage/reg_bank/reg_bank[73] , \iRF_stage/reg_bank/reg_bank[74] ,
         \iRF_stage/reg_bank/reg_bank[75] , \iRF_stage/reg_bank/reg_bank[76] ,
         \iRF_stage/reg_bank/reg_bank[77] , \iRF_stage/reg_bank/reg_bank[78] ,
         \iRF_stage/reg_bank/reg_bank[79] , \iRF_stage/reg_bank/reg_bank[80] ,
         \iRF_stage/reg_bank/reg_bank[81] , \iRF_stage/reg_bank/reg_bank[82] ,
         \iRF_stage/reg_bank/reg_bank[83] , \iRF_stage/reg_bank/reg_bank[84] ,
         \iRF_stage/reg_bank/reg_bank[85] , \iRF_stage/reg_bank/reg_bank[86] ,
         \iRF_stage/reg_bank/reg_bank[87] , \iRF_stage/reg_bank/reg_bank[88] ,
         \iRF_stage/reg_bank/reg_bank[89] , \iRF_stage/reg_bank/reg_bank[90] ,
         \iRF_stage/reg_bank/reg_bank[91] , \iRF_stage/reg_bank/reg_bank[92] ,
         \iRF_stage/reg_bank/reg_bank[93] , \iRF_stage/reg_bank/reg_bank[94] ,
         \iRF_stage/reg_bank/reg_bank[95] , \iRF_stage/reg_bank/reg_bank[96] ,
         \iRF_stage/reg_bank/reg_bank[97] , \iRF_stage/reg_bank/reg_bank[98] ,
         \iRF_stage/reg_bank/reg_bank[99] , \iRF_stage/reg_bank/reg_bank[100] ,
         \iRF_stage/reg_bank/reg_bank[101] ,
         \iRF_stage/reg_bank/reg_bank[102] ,
         \iRF_stage/reg_bank/reg_bank[103] ,
         \iRF_stage/reg_bank/reg_bank[104] ,
         \iRF_stage/reg_bank/reg_bank[105] ,
         \iRF_stage/reg_bank/reg_bank[106] ,
         \iRF_stage/reg_bank/reg_bank[107] ,
         \iRF_stage/reg_bank/reg_bank[108] ,
         \iRF_stage/reg_bank/reg_bank[109] ,
         \iRF_stage/reg_bank/reg_bank[110] ,
         \iRF_stage/reg_bank/reg_bank[111] ,
         \iRF_stage/reg_bank/reg_bank[112] ,
         \iRF_stage/reg_bank/reg_bank[113] ,
         \iRF_stage/reg_bank/reg_bank[114] ,
         \iRF_stage/reg_bank/reg_bank[115] ,
         \iRF_stage/reg_bank/reg_bank[116] ,
         \iRF_stage/reg_bank/reg_bank[117] ,
         \iRF_stage/reg_bank/reg_bank[118] ,
         \iRF_stage/reg_bank/reg_bank[119] ,
         \iRF_stage/reg_bank/reg_bank[120] ,
         \iRF_stage/reg_bank/reg_bank[121] ,
         \iRF_stage/reg_bank/reg_bank[122] ,
         \iRF_stage/reg_bank/reg_bank[123] ,
         \iRF_stage/reg_bank/reg_bank[124] ,
         \iRF_stage/reg_bank/reg_bank[125] ,
         \iRF_stage/reg_bank/reg_bank[126] ,
         \iRF_stage/reg_bank/reg_bank[127] ,
         \iRF_stage/reg_bank/reg_bank[128] ,
         \iRF_stage/reg_bank/reg_bank[129] ,
         \iRF_stage/reg_bank/reg_bank[130] ,
         \iRF_stage/reg_bank/reg_bank[131] ,
         \iRF_stage/reg_bank/reg_bank[132] ,
         \iRF_stage/reg_bank/reg_bank[133] ,
         \iRF_stage/reg_bank/reg_bank[134] ,
         \iRF_stage/reg_bank/reg_bank[135] ,
         \iRF_stage/reg_bank/reg_bank[136] ,
         \iRF_stage/reg_bank/reg_bank[137] ,
         \iRF_stage/reg_bank/reg_bank[138] ,
         \iRF_stage/reg_bank/reg_bank[139] ,
         \iRF_stage/reg_bank/reg_bank[140] ,
         \iRF_stage/reg_bank/reg_bank[141] ,
         \iRF_stage/reg_bank/reg_bank[142] ,
         \iRF_stage/reg_bank/reg_bank[143] ,
         \iRF_stage/reg_bank/reg_bank[144] ,
         \iRF_stage/reg_bank/reg_bank[145] ,
         \iRF_stage/reg_bank/reg_bank[146] ,
         \iRF_stage/reg_bank/reg_bank[147] ,
         \iRF_stage/reg_bank/reg_bank[148] ,
         \iRF_stage/reg_bank/reg_bank[149] ,
         \iRF_stage/reg_bank/reg_bank[150] ,
         \iRF_stage/reg_bank/reg_bank[151] ,
         \iRF_stage/reg_bank/reg_bank[152] ,
         \iRF_stage/reg_bank/reg_bank[153] ,
         \iRF_stage/reg_bank/reg_bank[154] ,
         \iRF_stage/reg_bank/reg_bank[155] ,
         \iRF_stage/reg_bank/reg_bank[156] ,
         \iRF_stage/reg_bank/reg_bank[157] ,
         \iRF_stage/reg_bank/reg_bank[158] ,
         \iRF_stage/reg_bank/reg_bank[159] ,
         \iRF_stage/reg_bank/reg_bank[160] ,
         \iRF_stage/reg_bank/reg_bank[161] ,
         \iRF_stage/reg_bank/reg_bank[162] ,
         \iRF_stage/reg_bank/reg_bank[163] ,
         \iRF_stage/reg_bank/reg_bank[164] ,
         \iRF_stage/reg_bank/reg_bank[165] ,
         \iRF_stage/reg_bank/reg_bank[166] ,
         \iRF_stage/reg_bank/reg_bank[167] ,
         \iRF_stage/reg_bank/reg_bank[168] ,
         \iRF_stage/reg_bank/reg_bank[169] ,
         \iRF_stage/reg_bank/reg_bank[170] ,
         \iRF_stage/reg_bank/reg_bank[171] ,
         \iRF_stage/reg_bank/reg_bank[172] ,
         \iRF_stage/reg_bank/reg_bank[173] ,
         \iRF_stage/reg_bank/reg_bank[174] ,
         \iRF_stage/reg_bank/reg_bank[175] ,
         \iRF_stage/reg_bank/reg_bank[176] ,
         \iRF_stage/reg_bank/reg_bank[177] ,
         \iRF_stage/reg_bank/reg_bank[178] ,
         \iRF_stage/reg_bank/reg_bank[179] ,
         \iRF_stage/reg_bank/reg_bank[180] ,
         \iRF_stage/reg_bank/reg_bank[181] ,
         \iRF_stage/reg_bank/reg_bank[182] ,
         \iRF_stage/reg_bank/reg_bank[183] ,
         \iRF_stage/reg_bank/reg_bank[184] ,
         \iRF_stage/reg_bank/reg_bank[185] ,
         \iRF_stage/reg_bank/reg_bank[186] ,
         \iRF_stage/reg_bank/reg_bank[187] ,
         \iRF_stage/reg_bank/reg_bank[188] ,
         \iRF_stage/reg_bank/reg_bank[189] ,
         \iRF_stage/reg_bank/reg_bank[190] ,
         \iRF_stage/reg_bank/reg_bank[191] ,
         \iRF_stage/reg_bank/reg_bank[192] ,
         \iRF_stage/reg_bank/reg_bank[193] ,
         \iRF_stage/reg_bank/reg_bank[194] ,
         \iRF_stage/reg_bank/reg_bank[195] ,
         \iRF_stage/reg_bank/reg_bank[196] ,
         \iRF_stage/reg_bank/reg_bank[197] ,
         \iRF_stage/reg_bank/reg_bank[198] ,
         \iRF_stage/reg_bank/reg_bank[199] ,
         \iRF_stage/reg_bank/reg_bank[200] ,
         \iRF_stage/reg_bank/reg_bank[201] ,
         \iRF_stage/reg_bank/reg_bank[202] ,
         \iRF_stage/reg_bank/reg_bank[203] ,
         \iRF_stage/reg_bank/reg_bank[204] ,
         \iRF_stage/reg_bank/reg_bank[205] ,
         \iRF_stage/reg_bank/reg_bank[206] ,
         \iRF_stage/reg_bank/reg_bank[207] ,
         \iRF_stage/reg_bank/reg_bank[208] ,
         \iRF_stage/reg_bank/reg_bank[209] ,
         \iRF_stage/reg_bank/reg_bank[210] ,
         \iRF_stage/reg_bank/reg_bank[211] ,
         \iRF_stage/reg_bank/reg_bank[212] ,
         \iRF_stage/reg_bank/reg_bank[213] ,
         \iRF_stage/reg_bank/reg_bank[214] ,
         \iRF_stage/reg_bank/reg_bank[215] ,
         \iRF_stage/reg_bank/reg_bank[216] ,
         \iRF_stage/reg_bank/reg_bank[217] ,
         \iRF_stage/reg_bank/reg_bank[218] ,
         \iRF_stage/reg_bank/reg_bank[219] ,
         \iRF_stage/reg_bank/reg_bank[220] ,
         \iRF_stage/reg_bank/reg_bank[221] ,
         \iRF_stage/reg_bank/reg_bank[222] ,
         \iRF_stage/reg_bank/reg_bank[223] ,
         \iRF_stage/reg_bank/reg_bank[224] ,
         \iRF_stage/reg_bank/reg_bank[225] ,
         \iRF_stage/reg_bank/reg_bank[226] ,
         \iRF_stage/reg_bank/reg_bank[227] ,
         \iRF_stage/reg_bank/reg_bank[228] ,
         \iRF_stage/reg_bank/reg_bank[229] ,
         \iRF_stage/reg_bank/reg_bank[230] ,
         \iRF_stage/reg_bank/reg_bank[231] ,
         \iRF_stage/reg_bank/reg_bank[232] ,
         \iRF_stage/reg_bank/reg_bank[233] ,
         \iRF_stage/reg_bank/reg_bank[234] ,
         \iRF_stage/reg_bank/reg_bank[235] ,
         \iRF_stage/reg_bank/reg_bank[236] ,
         \iRF_stage/reg_bank/reg_bank[237] ,
         \iRF_stage/reg_bank/reg_bank[238] ,
         \iRF_stage/reg_bank/reg_bank[239] ,
         \iRF_stage/reg_bank/reg_bank[240] ,
         \iRF_stage/reg_bank/reg_bank[241] ,
         \iRF_stage/reg_bank/reg_bank[242] ,
         \iRF_stage/reg_bank/reg_bank[243] ,
         \iRF_stage/reg_bank/reg_bank[244] ,
         \iRF_stage/reg_bank/reg_bank[245] ,
         \iRF_stage/reg_bank/reg_bank[246] ,
         \iRF_stage/reg_bank/reg_bank[247] ,
         \iRF_stage/reg_bank/reg_bank[248] ,
         \iRF_stage/reg_bank/reg_bank[249] ,
         \iRF_stage/reg_bank/reg_bank[250] ,
         \iRF_stage/reg_bank/reg_bank[251] ,
         \iRF_stage/reg_bank/reg_bank[252] ,
         \iRF_stage/reg_bank/reg_bank[253] ,
         \iRF_stage/reg_bank/reg_bank[254] ,
         \iRF_stage/reg_bank/reg_bank[255] ,
         \iRF_stage/reg_bank/reg_bank[256] ,
         \iRF_stage/reg_bank/reg_bank[257] ,
         \iRF_stage/reg_bank/reg_bank[258] ,
         \iRF_stage/reg_bank/reg_bank[259] ,
         \iRF_stage/reg_bank/reg_bank[260] ,
         \iRF_stage/reg_bank/reg_bank[261] ,
         \iRF_stage/reg_bank/reg_bank[262] ,
         \iRF_stage/reg_bank/reg_bank[263] ,
         \iRF_stage/reg_bank/reg_bank[264] ,
         \iRF_stage/reg_bank/reg_bank[265] ,
         \iRF_stage/reg_bank/reg_bank[266] ,
         \iRF_stage/reg_bank/reg_bank[267] ,
         \iRF_stage/reg_bank/reg_bank[268] ,
         \iRF_stage/reg_bank/reg_bank[269] ,
         \iRF_stage/reg_bank/reg_bank[270] ,
         \iRF_stage/reg_bank/reg_bank[271] ,
         \iRF_stage/reg_bank/reg_bank[272] ,
         \iRF_stage/reg_bank/reg_bank[273] ,
         \iRF_stage/reg_bank/reg_bank[274] ,
         \iRF_stage/reg_bank/reg_bank[275] ,
         \iRF_stage/reg_bank/reg_bank[276] ,
         \iRF_stage/reg_bank/reg_bank[277] ,
         \iRF_stage/reg_bank/reg_bank[278] ,
         \iRF_stage/reg_bank/reg_bank[279] ,
         \iRF_stage/reg_bank/reg_bank[280] ,
         \iRF_stage/reg_bank/reg_bank[281] ,
         \iRF_stage/reg_bank/reg_bank[282] ,
         \iRF_stage/reg_bank/reg_bank[283] ,
         \iRF_stage/reg_bank/reg_bank[284] ,
         \iRF_stage/reg_bank/reg_bank[285] ,
         \iRF_stage/reg_bank/reg_bank[286] ,
         \iRF_stage/reg_bank/reg_bank[287] ,
         \iRF_stage/reg_bank/reg_bank[288] ,
         \iRF_stage/reg_bank/reg_bank[289] ,
         \iRF_stage/reg_bank/reg_bank[290] ,
         \iRF_stage/reg_bank/reg_bank[291] ,
         \iRF_stage/reg_bank/reg_bank[292] ,
         \iRF_stage/reg_bank/reg_bank[293] ,
         \iRF_stage/reg_bank/reg_bank[294] ,
         \iRF_stage/reg_bank/reg_bank[295] ,
         \iRF_stage/reg_bank/reg_bank[296] ,
         \iRF_stage/reg_bank/reg_bank[297] ,
         \iRF_stage/reg_bank/reg_bank[298] ,
         \iRF_stage/reg_bank/reg_bank[299] ,
         \iRF_stage/reg_bank/reg_bank[300] ,
         \iRF_stage/reg_bank/reg_bank[301] ,
         \iRF_stage/reg_bank/reg_bank[302] ,
         \iRF_stage/reg_bank/reg_bank[303] ,
         \iRF_stage/reg_bank/reg_bank[304] ,
         \iRF_stage/reg_bank/reg_bank[305] ,
         \iRF_stage/reg_bank/reg_bank[306] ,
         \iRF_stage/reg_bank/reg_bank[307] ,
         \iRF_stage/reg_bank/reg_bank[308] ,
         \iRF_stage/reg_bank/reg_bank[309] ,
         \iRF_stage/reg_bank/reg_bank[310] ,
         \iRF_stage/reg_bank/reg_bank[311] ,
         \iRF_stage/reg_bank/reg_bank[312] ,
         \iRF_stage/reg_bank/reg_bank[313] ,
         \iRF_stage/reg_bank/reg_bank[314] ,
         \iRF_stage/reg_bank/reg_bank[315] ,
         \iRF_stage/reg_bank/reg_bank[316] ,
         \iRF_stage/reg_bank/reg_bank[317] ,
         \iRF_stage/reg_bank/reg_bank[318] ,
         \iRF_stage/reg_bank/reg_bank[319] ,
         \iRF_stage/reg_bank/reg_bank[320] ,
         \iRF_stage/reg_bank/reg_bank[321] ,
         \iRF_stage/reg_bank/reg_bank[322] ,
         \iRF_stage/reg_bank/reg_bank[323] ,
         \iRF_stage/reg_bank/reg_bank[324] ,
         \iRF_stage/reg_bank/reg_bank[325] ,
         \iRF_stage/reg_bank/reg_bank[326] ,
         \iRF_stage/reg_bank/reg_bank[327] ,
         \iRF_stage/reg_bank/reg_bank[328] ,
         \iRF_stage/reg_bank/reg_bank[329] ,
         \iRF_stage/reg_bank/reg_bank[330] ,
         \iRF_stage/reg_bank/reg_bank[331] ,
         \iRF_stage/reg_bank/reg_bank[332] ,
         \iRF_stage/reg_bank/reg_bank[333] ,
         \iRF_stage/reg_bank/reg_bank[334] ,
         \iRF_stage/reg_bank/reg_bank[335] ,
         \iRF_stage/reg_bank/reg_bank[336] ,
         \iRF_stage/reg_bank/reg_bank[337] ,
         \iRF_stage/reg_bank/reg_bank[338] ,
         \iRF_stage/reg_bank/reg_bank[339] ,
         \iRF_stage/reg_bank/reg_bank[340] ,
         \iRF_stage/reg_bank/reg_bank[341] ,
         \iRF_stage/reg_bank/reg_bank[342] ,
         \iRF_stage/reg_bank/reg_bank[343] ,
         \iRF_stage/reg_bank/reg_bank[344] ,
         \iRF_stage/reg_bank/reg_bank[345] ,
         \iRF_stage/reg_bank/reg_bank[346] ,
         \iRF_stage/reg_bank/reg_bank[347] ,
         \iRF_stage/reg_bank/reg_bank[348] ,
         \iRF_stage/reg_bank/reg_bank[349] ,
         \iRF_stage/reg_bank/reg_bank[350] ,
         \iRF_stage/reg_bank/reg_bank[351] ,
         \iRF_stage/reg_bank/reg_bank[352] ,
         \iRF_stage/reg_bank/reg_bank[353] ,
         \iRF_stage/reg_bank/reg_bank[354] ,
         \iRF_stage/reg_bank/reg_bank[355] ,
         \iRF_stage/reg_bank/reg_bank[356] ,
         \iRF_stage/reg_bank/reg_bank[357] ,
         \iRF_stage/reg_bank/reg_bank[358] ,
         \iRF_stage/reg_bank/reg_bank[359] ,
         \iRF_stage/reg_bank/reg_bank[360] ,
         \iRF_stage/reg_bank/reg_bank[361] ,
         \iRF_stage/reg_bank/reg_bank[362] ,
         \iRF_stage/reg_bank/reg_bank[363] ,
         \iRF_stage/reg_bank/reg_bank[364] ,
         \iRF_stage/reg_bank/reg_bank[365] ,
         \iRF_stage/reg_bank/reg_bank[366] ,
         \iRF_stage/reg_bank/reg_bank[367] ,
         \iRF_stage/reg_bank/reg_bank[368] ,
         \iRF_stage/reg_bank/reg_bank[369] ,
         \iRF_stage/reg_bank/reg_bank[370] ,
         \iRF_stage/reg_bank/reg_bank[371] ,
         \iRF_stage/reg_bank/reg_bank[372] ,
         \iRF_stage/reg_bank/reg_bank[373] ,
         \iRF_stage/reg_bank/reg_bank[374] ,
         \iRF_stage/reg_bank/reg_bank[375] ,
         \iRF_stage/reg_bank/reg_bank[376] ,
         \iRF_stage/reg_bank/reg_bank[377] ,
         \iRF_stage/reg_bank/reg_bank[378] ,
         \iRF_stage/reg_bank/reg_bank[379] ,
         \iRF_stage/reg_bank/reg_bank[380] ,
         \iRF_stage/reg_bank/reg_bank[381] ,
         \iRF_stage/reg_bank/reg_bank[382] ,
         \iRF_stage/reg_bank/reg_bank[383] ,
         \iRF_stage/reg_bank/reg_bank[384] ,
         \iRF_stage/reg_bank/reg_bank[385] ,
         \iRF_stage/reg_bank/reg_bank[386] ,
         \iRF_stage/reg_bank/reg_bank[387] ,
         \iRF_stage/reg_bank/reg_bank[388] ,
         \iRF_stage/reg_bank/reg_bank[389] ,
         \iRF_stage/reg_bank/reg_bank[390] ,
         \iRF_stage/reg_bank/reg_bank[391] ,
         \iRF_stage/reg_bank/reg_bank[392] ,
         \iRF_stage/reg_bank/reg_bank[393] ,
         \iRF_stage/reg_bank/reg_bank[394] ,
         \iRF_stage/reg_bank/reg_bank[395] ,
         \iRF_stage/reg_bank/reg_bank[396] ,
         \iRF_stage/reg_bank/reg_bank[397] ,
         \iRF_stage/reg_bank/reg_bank[398] ,
         \iRF_stage/reg_bank/reg_bank[399] ,
         \iRF_stage/reg_bank/reg_bank[400] ,
         \iRF_stage/reg_bank/reg_bank[401] ,
         \iRF_stage/reg_bank/reg_bank[402] ,
         \iRF_stage/reg_bank/reg_bank[403] ,
         \iRF_stage/reg_bank/reg_bank[404] ,
         \iRF_stage/reg_bank/reg_bank[405] ,
         \iRF_stage/reg_bank/reg_bank[406] ,
         \iRF_stage/reg_bank/reg_bank[407] ,
         \iRF_stage/reg_bank/reg_bank[408] ,
         \iRF_stage/reg_bank/reg_bank[409] ,
         \iRF_stage/reg_bank/reg_bank[410] ,
         \iRF_stage/reg_bank/reg_bank[411] ,
         \iRF_stage/reg_bank/reg_bank[412] ,
         \iRF_stage/reg_bank/reg_bank[413] ,
         \iRF_stage/reg_bank/reg_bank[414] ,
         \iRF_stage/reg_bank/reg_bank[415] ,
         \iRF_stage/reg_bank/reg_bank[416] ,
         \iRF_stage/reg_bank/reg_bank[417] ,
         \iRF_stage/reg_bank/reg_bank[418] ,
         \iRF_stage/reg_bank/reg_bank[419] ,
         \iRF_stage/reg_bank/reg_bank[420] ,
         \iRF_stage/reg_bank/reg_bank[421] ,
         \iRF_stage/reg_bank/reg_bank[422] ,
         \iRF_stage/reg_bank/reg_bank[423] ,
         \iRF_stage/reg_bank/reg_bank[424] ,
         \iRF_stage/reg_bank/reg_bank[425] ,
         \iRF_stage/reg_bank/reg_bank[426] ,
         \iRF_stage/reg_bank/reg_bank[427] ,
         \iRF_stage/reg_bank/reg_bank[428] ,
         \iRF_stage/reg_bank/reg_bank[429] ,
         \iRF_stage/reg_bank/reg_bank[430] ,
         \iRF_stage/reg_bank/reg_bank[431] ,
         \iRF_stage/reg_bank/reg_bank[432] ,
         \iRF_stage/reg_bank/reg_bank[433] ,
         \iRF_stage/reg_bank/reg_bank[434] ,
         \iRF_stage/reg_bank/reg_bank[435] ,
         \iRF_stage/reg_bank/reg_bank[436] ,
         \iRF_stage/reg_bank/reg_bank[437] ,
         \iRF_stage/reg_bank/reg_bank[438] ,
         \iRF_stage/reg_bank/reg_bank[439] ,
         \iRF_stage/reg_bank/reg_bank[440] ,
         \iRF_stage/reg_bank/reg_bank[441] ,
         \iRF_stage/reg_bank/reg_bank[442] ,
         \iRF_stage/reg_bank/reg_bank[443] ,
         \iRF_stage/reg_bank/reg_bank[444] ,
         \iRF_stage/reg_bank/reg_bank[445] ,
         \iRF_stage/reg_bank/reg_bank[446] ,
         \iRF_stage/reg_bank/reg_bank[447] ,
         \iRF_stage/reg_bank/reg_bank[448] ,
         \iRF_stage/reg_bank/reg_bank[449] ,
         \iRF_stage/reg_bank/reg_bank[450] ,
         \iRF_stage/reg_bank/reg_bank[451] ,
         \iRF_stage/reg_bank/reg_bank[452] ,
         \iRF_stage/reg_bank/reg_bank[453] ,
         \iRF_stage/reg_bank/reg_bank[454] ,
         \iRF_stage/reg_bank/reg_bank[455] ,
         \iRF_stage/reg_bank/reg_bank[456] ,
         \iRF_stage/reg_bank/reg_bank[457] ,
         \iRF_stage/reg_bank/reg_bank[458] ,
         \iRF_stage/reg_bank/reg_bank[459] ,
         \iRF_stage/reg_bank/reg_bank[460] ,
         \iRF_stage/reg_bank/reg_bank[461] ,
         \iRF_stage/reg_bank/reg_bank[462] ,
         \iRF_stage/reg_bank/reg_bank[463] ,
         \iRF_stage/reg_bank/reg_bank[464] ,
         \iRF_stage/reg_bank/reg_bank[465] ,
         \iRF_stage/reg_bank/reg_bank[466] ,
         \iRF_stage/reg_bank/reg_bank[467] ,
         \iRF_stage/reg_bank/reg_bank[468] ,
         \iRF_stage/reg_bank/reg_bank[469] ,
         \iRF_stage/reg_bank/reg_bank[470] ,
         \iRF_stage/reg_bank/reg_bank[471] ,
         \iRF_stage/reg_bank/reg_bank[472] ,
         \iRF_stage/reg_bank/reg_bank[473] ,
         \iRF_stage/reg_bank/reg_bank[474] ,
         \iRF_stage/reg_bank/reg_bank[475] ,
         \iRF_stage/reg_bank/reg_bank[476] ,
         \iRF_stage/reg_bank/reg_bank[477] ,
         \iRF_stage/reg_bank/reg_bank[478] ,
         \iRF_stage/reg_bank/reg_bank[479] ,
         \iRF_stage/reg_bank/reg_bank[480] ,
         \iRF_stage/reg_bank/reg_bank[481] ,
         \iRF_stage/reg_bank/reg_bank[482] ,
         \iRF_stage/reg_bank/reg_bank[483] ,
         \iRF_stage/reg_bank/reg_bank[484] ,
         \iRF_stage/reg_bank/reg_bank[485] ,
         \iRF_stage/reg_bank/reg_bank[486] ,
         \iRF_stage/reg_bank/reg_bank[487] ,
         \iRF_stage/reg_bank/reg_bank[488] ,
         \iRF_stage/reg_bank/reg_bank[489] ,
         \iRF_stage/reg_bank/reg_bank[490] ,
         \iRF_stage/reg_bank/reg_bank[491] ,
         \iRF_stage/reg_bank/reg_bank[492] ,
         \iRF_stage/reg_bank/reg_bank[493] ,
         \iRF_stage/reg_bank/reg_bank[494] ,
         \iRF_stage/reg_bank/reg_bank[495] ,
         \iRF_stage/reg_bank/reg_bank[496] ,
         \iRF_stage/reg_bank/reg_bank[497] ,
         \iRF_stage/reg_bank/reg_bank[498] ,
         \iRF_stage/reg_bank/reg_bank[499] ,
         \iRF_stage/reg_bank/reg_bank[500] ,
         \iRF_stage/reg_bank/reg_bank[501] ,
         \iRF_stage/reg_bank/reg_bank[502] ,
         \iRF_stage/reg_bank/reg_bank[503] ,
         \iRF_stage/reg_bank/reg_bank[504] ,
         \iRF_stage/reg_bank/reg_bank[505] ,
         \iRF_stage/reg_bank/reg_bank[506] ,
         \iRF_stage/reg_bank/reg_bank[507] ,
         \iRF_stage/reg_bank/reg_bank[508] ,
         \iRF_stage/reg_bank/reg_bank[509] ,
         \iRF_stage/reg_bank/reg_bank[510] ,
         \iRF_stage/reg_bank/reg_bank[511] ,
         \iRF_stage/reg_bank/reg_bank[512] ,
         \iRF_stage/reg_bank/reg_bank[513] ,
         \iRF_stage/reg_bank/reg_bank[514] ,
         \iRF_stage/reg_bank/reg_bank[515] ,
         \iRF_stage/reg_bank/reg_bank[516] ,
         \iRF_stage/reg_bank/reg_bank[517] ,
         \iRF_stage/reg_bank/reg_bank[518] ,
         \iRF_stage/reg_bank/reg_bank[519] ,
         \iRF_stage/reg_bank/reg_bank[520] ,
         \iRF_stage/reg_bank/reg_bank[521] ,
         \iRF_stage/reg_bank/reg_bank[522] ,
         \iRF_stage/reg_bank/reg_bank[523] ,
         \iRF_stage/reg_bank/reg_bank[524] ,
         \iRF_stage/reg_bank/reg_bank[525] ,
         \iRF_stage/reg_bank/reg_bank[526] ,
         \iRF_stage/reg_bank/reg_bank[527] ,
         \iRF_stage/reg_bank/reg_bank[528] ,
         \iRF_stage/reg_bank/reg_bank[529] ,
         \iRF_stage/reg_bank/reg_bank[530] ,
         \iRF_stage/reg_bank/reg_bank[531] ,
         \iRF_stage/reg_bank/reg_bank[532] ,
         \iRF_stage/reg_bank/reg_bank[533] ,
         \iRF_stage/reg_bank/reg_bank[534] ,
         \iRF_stage/reg_bank/reg_bank[535] ,
         \iRF_stage/reg_bank/reg_bank[536] ,
         \iRF_stage/reg_bank/reg_bank[537] ,
         \iRF_stage/reg_bank/reg_bank[538] ,
         \iRF_stage/reg_bank/reg_bank[539] ,
         \iRF_stage/reg_bank/reg_bank[540] ,
         \iRF_stage/reg_bank/reg_bank[541] ,
         \iRF_stage/reg_bank/reg_bank[542] ,
         \iRF_stage/reg_bank/reg_bank[543] ,
         \iRF_stage/reg_bank/reg_bank[544] ,
         \iRF_stage/reg_bank/reg_bank[545] ,
         \iRF_stage/reg_bank/reg_bank[546] ,
         \iRF_stage/reg_bank/reg_bank[547] ,
         \iRF_stage/reg_bank/reg_bank[548] ,
         \iRF_stage/reg_bank/reg_bank[549] ,
         \iRF_stage/reg_bank/reg_bank[550] ,
         \iRF_stage/reg_bank/reg_bank[551] ,
         \iRF_stage/reg_bank/reg_bank[552] ,
         \iRF_stage/reg_bank/reg_bank[553] ,
         \iRF_stage/reg_bank/reg_bank[554] ,
         \iRF_stage/reg_bank/reg_bank[555] ,
         \iRF_stage/reg_bank/reg_bank[556] ,
         \iRF_stage/reg_bank/reg_bank[557] ,
         \iRF_stage/reg_bank/reg_bank[558] ,
         \iRF_stage/reg_bank/reg_bank[559] ,
         \iRF_stage/reg_bank/reg_bank[560] ,
         \iRF_stage/reg_bank/reg_bank[561] ,
         \iRF_stage/reg_bank/reg_bank[562] ,
         \iRF_stage/reg_bank/reg_bank[563] ,
         \iRF_stage/reg_bank/reg_bank[564] ,
         \iRF_stage/reg_bank/reg_bank[565] ,
         \iRF_stage/reg_bank/reg_bank[566] ,
         \iRF_stage/reg_bank/reg_bank[567] ,
         \iRF_stage/reg_bank/reg_bank[568] ,
         \iRF_stage/reg_bank/reg_bank[569] ,
         \iRF_stage/reg_bank/reg_bank[570] ,
         \iRF_stage/reg_bank/reg_bank[571] ,
         \iRF_stage/reg_bank/reg_bank[572] ,
         \iRF_stage/reg_bank/reg_bank[573] ,
         \iRF_stage/reg_bank/reg_bank[574] ,
         \iRF_stage/reg_bank/reg_bank[575] ,
         \iRF_stage/reg_bank/reg_bank[576] ,
         \iRF_stage/reg_bank/reg_bank[577] ,
         \iRF_stage/reg_bank/reg_bank[578] ,
         \iRF_stage/reg_bank/reg_bank[579] ,
         \iRF_stage/reg_bank/reg_bank[580] ,
         \iRF_stage/reg_bank/reg_bank[581] ,
         \iRF_stage/reg_bank/reg_bank[582] ,
         \iRF_stage/reg_bank/reg_bank[583] ,
         \iRF_stage/reg_bank/reg_bank[584] ,
         \iRF_stage/reg_bank/reg_bank[585] ,
         \iRF_stage/reg_bank/reg_bank[586] ,
         \iRF_stage/reg_bank/reg_bank[587] ,
         \iRF_stage/reg_bank/reg_bank[588] ,
         \iRF_stage/reg_bank/reg_bank[589] ,
         \iRF_stage/reg_bank/reg_bank[590] ,
         \iRF_stage/reg_bank/reg_bank[591] ,
         \iRF_stage/reg_bank/reg_bank[592] ,
         \iRF_stage/reg_bank/reg_bank[593] ,
         \iRF_stage/reg_bank/reg_bank[594] ,
         \iRF_stage/reg_bank/reg_bank[595] ,
         \iRF_stage/reg_bank/reg_bank[596] ,
         \iRF_stage/reg_bank/reg_bank[597] ,
         \iRF_stage/reg_bank/reg_bank[598] ,
         \iRF_stage/reg_bank/reg_bank[599] ,
         \iRF_stage/reg_bank/reg_bank[600] ,
         \iRF_stage/reg_bank/reg_bank[601] ,
         \iRF_stage/reg_bank/reg_bank[602] ,
         \iRF_stage/reg_bank/reg_bank[603] ,
         \iRF_stage/reg_bank/reg_bank[604] ,
         \iRF_stage/reg_bank/reg_bank[605] ,
         \iRF_stage/reg_bank/reg_bank[606] ,
         \iRF_stage/reg_bank/reg_bank[607] ,
         \iRF_stage/reg_bank/reg_bank[608] ,
         \iRF_stage/reg_bank/reg_bank[609] ,
         \iRF_stage/reg_bank/reg_bank[610] ,
         \iRF_stage/reg_bank/reg_bank[611] ,
         \iRF_stage/reg_bank/reg_bank[612] ,
         \iRF_stage/reg_bank/reg_bank[613] ,
         \iRF_stage/reg_bank/reg_bank[614] ,
         \iRF_stage/reg_bank/reg_bank[615] ,
         \iRF_stage/reg_bank/reg_bank[616] ,
         \iRF_stage/reg_bank/reg_bank[617] ,
         \iRF_stage/reg_bank/reg_bank[618] ,
         \iRF_stage/reg_bank/reg_bank[619] ,
         \iRF_stage/reg_bank/reg_bank[620] ,
         \iRF_stage/reg_bank/reg_bank[621] ,
         \iRF_stage/reg_bank/reg_bank[622] ,
         \iRF_stage/reg_bank/reg_bank[623] ,
         \iRF_stage/reg_bank/reg_bank[624] ,
         \iRF_stage/reg_bank/reg_bank[625] ,
         \iRF_stage/reg_bank/reg_bank[626] ,
         \iRF_stage/reg_bank/reg_bank[627] ,
         \iRF_stage/reg_bank/reg_bank[628] ,
         \iRF_stage/reg_bank/reg_bank[629] ,
         \iRF_stage/reg_bank/reg_bank[630] ,
         \iRF_stage/reg_bank/reg_bank[631] ,
         \iRF_stage/reg_bank/reg_bank[632] ,
         \iRF_stage/reg_bank/reg_bank[633] ,
         \iRF_stage/reg_bank/reg_bank[634] ,
         \iRF_stage/reg_bank/reg_bank[635] ,
         \iRF_stage/reg_bank/reg_bank[636] ,
         \iRF_stage/reg_bank/reg_bank[637] ,
         \iRF_stage/reg_bank/reg_bank[638] ,
         \iRF_stage/reg_bank/reg_bank[639] ,
         \iRF_stage/reg_bank/reg_bank[640] ,
         \iRF_stage/reg_bank/reg_bank[641] ,
         \iRF_stage/reg_bank/reg_bank[642] ,
         \iRF_stage/reg_bank/reg_bank[643] ,
         \iRF_stage/reg_bank/reg_bank[644] ,
         \iRF_stage/reg_bank/reg_bank[645] ,
         \iRF_stage/reg_bank/reg_bank[646] ,
         \iRF_stage/reg_bank/reg_bank[647] ,
         \iRF_stage/reg_bank/reg_bank[648] ,
         \iRF_stage/reg_bank/reg_bank[649] ,
         \iRF_stage/reg_bank/reg_bank[650] ,
         \iRF_stage/reg_bank/reg_bank[651] ,
         \iRF_stage/reg_bank/reg_bank[652] ,
         \iRF_stage/reg_bank/reg_bank[653] ,
         \iRF_stage/reg_bank/reg_bank[654] ,
         \iRF_stage/reg_bank/reg_bank[655] ,
         \iRF_stage/reg_bank/reg_bank[656] ,
         \iRF_stage/reg_bank/reg_bank[657] ,
         \iRF_stage/reg_bank/reg_bank[658] ,
         \iRF_stage/reg_bank/reg_bank[659] ,
         \iRF_stage/reg_bank/reg_bank[660] ,
         \iRF_stage/reg_bank/reg_bank[661] ,
         \iRF_stage/reg_bank/reg_bank[662] ,
         \iRF_stage/reg_bank/reg_bank[663] ,
         \iRF_stage/reg_bank/reg_bank[664] ,
         \iRF_stage/reg_bank/reg_bank[665] ,
         \iRF_stage/reg_bank/reg_bank[666] ,
         \iRF_stage/reg_bank/reg_bank[667] ,
         \iRF_stage/reg_bank/reg_bank[668] ,
         \iRF_stage/reg_bank/reg_bank[669] ,
         \iRF_stage/reg_bank/reg_bank[670] ,
         \iRF_stage/reg_bank/reg_bank[671] ,
         \iRF_stage/reg_bank/reg_bank[672] ,
         \iRF_stage/reg_bank/reg_bank[673] ,
         \iRF_stage/reg_bank/reg_bank[674] ,
         \iRF_stage/reg_bank/reg_bank[675] ,
         \iRF_stage/reg_bank/reg_bank[676] ,
         \iRF_stage/reg_bank/reg_bank[677] ,
         \iRF_stage/reg_bank/reg_bank[678] ,
         \iRF_stage/reg_bank/reg_bank[679] ,
         \iRF_stage/reg_bank/reg_bank[680] ,
         \iRF_stage/reg_bank/reg_bank[681] ,
         \iRF_stage/reg_bank/reg_bank[682] ,
         \iRF_stage/reg_bank/reg_bank[683] ,
         \iRF_stage/reg_bank/reg_bank[684] ,
         \iRF_stage/reg_bank/reg_bank[685] ,
         \iRF_stage/reg_bank/reg_bank[686] ,
         \iRF_stage/reg_bank/reg_bank[687] ,
         \iRF_stage/reg_bank/reg_bank[688] ,
         \iRF_stage/reg_bank/reg_bank[689] ,
         \iRF_stage/reg_bank/reg_bank[690] ,
         \iRF_stage/reg_bank/reg_bank[691] ,
         \iRF_stage/reg_bank/reg_bank[692] ,
         \iRF_stage/reg_bank/reg_bank[693] ,
         \iRF_stage/reg_bank/reg_bank[694] ,
         \iRF_stage/reg_bank/reg_bank[695] ,
         \iRF_stage/reg_bank/reg_bank[696] ,
         \iRF_stage/reg_bank/reg_bank[697] ,
         \iRF_stage/reg_bank/reg_bank[698] ,
         \iRF_stage/reg_bank/reg_bank[699] ,
         \iRF_stage/reg_bank/reg_bank[700] ,
         \iRF_stage/reg_bank/reg_bank[701] ,
         \iRF_stage/reg_bank/reg_bank[702] ,
         \iRF_stage/reg_bank/reg_bank[703] ,
         \iRF_stage/reg_bank/reg_bank[704] ,
         \iRF_stage/reg_bank/reg_bank[705] ,
         \iRF_stage/reg_bank/reg_bank[706] ,
         \iRF_stage/reg_bank/reg_bank[707] ,
         \iRF_stage/reg_bank/reg_bank[708] ,
         \iRF_stage/reg_bank/reg_bank[709] ,
         \iRF_stage/reg_bank/reg_bank[710] ,
         \iRF_stage/reg_bank/reg_bank[711] ,
         \iRF_stage/reg_bank/reg_bank[712] ,
         \iRF_stage/reg_bank/reg_bank[713] ,
         \iRF_stage/reg_bank/reg_bank[714] ,
         \iRF_stage/reg_bank/reg_bank[715] ,
         \iRF_stage/reg_bank/reg_bank[716] ,
         \iRF_stage/reg_bank/reg_bank[717] ,
         \iRF_stage/reg_bank/reg_bank[718] ,
         \iRF_stage/reg_bank/reg_bank[719] ,
         \iRF_stage/reg_bank/reg_bank[720] ,
         \iRF_stage/reg_bank/reg_bank[721] ,
         \iRF_stage/reg_bank/reg_bank[722] ,
         \iRF_stage/reg_bank/reg_bank[723] ,
         \iRF_stage/reg_bank/reg_bank[724] ,
         \iRF_stage/reg_bank/reg_bank[725] ,
         \iRF_stage/reg_bank/reg_bank[726] ,
         \iRF_stage/reg_bank/reg_bank[727] ,
         \iRF_stage/reg_bank/reg_bank[728] ,
         \iRF_stage/reg_bank/reg_bank[729] ,
         \iRF_stage/reg_bank/reg_bank[730] ,
         \iRF_stage/reg_bank/reg_bank[731] ,
         \iRF_stage/reg_bank/reg_bank[732] ,
         \iRF_stage/reg_bank/reg_bank[733] ,
         \iRF_stage/reg_bank/reg_bank[734] ,
         \iRF_stage/reg_bank/reg_bank[735] ,
         \iRF_stage/reg_bank/reg_bank[736] ,
         \iRF_stage/reg_bank/reg_bank[737] ,
         \iRF_stage/reg_bank/reg_bank[738] ,
         \iRF_stage/reg_bank/reg_bank[739] ,
         \iRF_stage/reg_bank/reg_bank[740] ,
         \iRF_stage/reg_bank/reg_bank[741] ,
         \iRF_stage/reg_bank/reg_bank[742] ,
         \iRF_stage/reg_bank/reg_bank[743] ,
         \iRF_stage/reg_bank/reg_bank[744] ,
         \iRF_stage/reg_bank/reg_bank[745] ,
         \iRF_stage/reg_bank/reg_bank[746] ,
         \iRF_stage/reg_bank/reg_bank[747] ,
         \iRF_stage/reg_bank/reg_bank[748] ,
         \iRF_stage/reg_bank/reg_bank[749] ,
         \iRF_stage/reg_bank/reg_bank[750] ,
         \iRF_stage/reg_bank/reg_bank[751] ,
         \iRF_stage/reg_bank/reg_bank[752] ,
         \iRF_stage/reg_bank/reg_bank[753] ,
         \iRF_stage/reg_bank/reg_bank[754] ,
         \iRF_stage/reg_bank/reg_bank[755] ,
         \iRF_stage/reg_bank/reg_bank[756] ,
         \iRF_stage/reg_bank/reg_bank[757] ,
         \iRF_stage/reg_bank/reg_bank[758] ,
         \iRF_stage/reg_bank/reg_bank[759] ,
         \iRF_stage/reg_bank/reg_bank[760] ,
         \iRF_stage/reg_bank/reg_bank[761] ,
         \iRF_stage/reg_bank/reg_bank[762] ,
         \iRF_stage/reg_bank/reg_bank[763] ,
         \iRF_stage/reg_bank/reg_bank[764] ,
         \iRF_stage/reg_bank/reg_bank[765] ,
         \iRF_stage/reg_bank/reg_bank[766] ,
         \iRF_stage/reg_bank/reg_bank[767] ,
         \iRF_stage/reg_bank/reg_bank[768] ,
         \iRF_stage/reg_bank/reg_bank[769] ,
         \iRF_stage/reg_bank/reg_bank[770] ,
         \iRF_stage/reg_bank/reg_bank[771] ,
         \iRF_stage/reg_bank/reg_bank[772] ,
         \iRF_stage/reg_bank/reg_bank[773] ,
         \iRF_stage/reg_bank/reg_bank[774] ,
         \iRF_stage/reg_bank/reg_bank[775] ,
         \iRF_stage/reg_bank/reg_bank[776] ,
         \iRF_stage/reg_bank/reg_bank[777] ,
         \iRF_stage/reg_bank/reg_bank[778] ,
         \iRF_stage/reg_bank/reg_bank[779] ,
         \iRF_stage/reg_bank/reg_bank[780] ,
         \iRF_stage/reg_bank/reg_bank[781] ,
         \iRF_stage/reg_bank/reg_bank[782] ,
         \iRF_stage/reg_bank/reg_bank[783] ,
         \iRF_stage/reg_bank/reg_bank[784] ,
         \iRF_stage/reg_bank/reg_bank[785] ,
         \iRF_stage/reg_bank/reg_bank[786] ,
         \iRF_stage/reg_bank/reg_bank[787] ,
         \iRF_stage/reg_bank/reg_bank[788] ,
         \iRF_stage/reg_bank/reg_bank[789] ,
         \iRF_stage/reg_bank/reg_bank[790] ,
         \iRF_stage/reg_bank/reg_bank[791] ,
         \iRF_stage/reg_bank/reg_bank[792] ,
         \iRF_stage/reg_bank/reg_bank[793] ,
         \iRF_stage/reg_bank/reg_bank[794] ,
         \iRF_stage/reg_bank/reg_bank[795] ,
         \iRF_stage/reg_bank/reg_bank[796] ,
         \iRF_stage/reg_bank/reg_bank[797] ,
         \iRF_stage/reg_bank/reg_bank[798] ,
         \iRF_stage/reg_bank/reg_bank[799] ,
         \iRF_stage/reg_bank/reg_bank[800] ,
         \iRF_stage/reg_bank/reg_bank[801] ,
         \iRF_stage/reg_bank/reg_bank[802] ,
         \iRF_stage/reg_bank/reg_bank[803] ,
         \iRF_stage/reg_bank/reg_bank[804] ,
         \iRF_stage/reg_bank/reg_bank[805] ,
         \iRF_stage/reg_bank/reg_bank[806] ,
         \iRF_stage/reg_bank/reg_bank[807] ,
         \iRF_stage/reg_bank/reg_bank[808] ,
         \iRF_stage/reg_bank/reg_bank[809] ,
         \iRF_stage/reg_bank/reg_bank[810] ,
         \iRF_stage/reg_bank/reg_bank[811] ,
         \iRF_stage/reg_bank/reg_bank[812] ,
         \iRF_stage/reg_bank/reg_bank[813] ,
         \iRF_stage/reg_bank/reg_bank[814] ,
         \iRF_stage/reg_bank/reg_bank[815] ,
         \iRF_stage/reg_bank/reg_bank[816] ,
         \iRF_stage/reg_bank/reg_bank[817] ,
         \iRF_stage/reg_bank/reg_bank[818] ,
         \iRF_stage/reg_bank/reg_bank[819] ,
         \iRF_stage/reg_bank/reg_bank[820] ,
         \iRF_stage/reg_bank/reg_bank[821] ,
         \iRF_stage/reg_bank/reg_bank[822] ,
         \iRF_stage/reg_bank/reg_bank[823] ,
         \iRF_stage/reg_bank/reg_bank[824] ,
         \iRF_stage/reg_bank/reg_bank[825] ,
         \iRF_stage/reg_bank/reg_bank[826] ,
         \iRF_stage/reg_bank/reg_bank[827] ,
         \iRF_stage/reg_bank/reg_bank[828] ,
         \iRF_stage/reg_bank/reg_bank[829] ,
         \iRF_stage/reg_bank/reg_bank[830] ,
         \iRF_stage/reg_bank/reg_bank[831] ,
         \iRF_stage/reg_bank/reg_bank[832] ,
         \iRF_stage/reg_bank/reg_bank[833] ,
         \iRF_stage/reg_bank/reg_bank[834] ,
         \iRF_stage/reg_bank/reg_bank[835] ,
         \iRF_stage/reg_bank/reg_bank[836] ,
         \iRF_stage/reg_bank/reg_bank[837] ,
         \iRF_stage/reg_bank/reg_bank[838] ,
         \iRF_stage/reg_bank/reg_bank[839] ,
         \iRF_stage/reg_bank/reg_bank[840] ,
         \iRF_stage/reg_bank/reg_bank[841] ,
         \iRF_stage/reg_bank/reg_bank[842] ,
         \iRF_stage/reg_bank/reg_bank[843] ,
         \iRF_stage/reg_bank/reg_bank[844] ,
         \iRF_stage/reg_bank/reg_bank[845] ,
         \iRF_stage/reg_bank/reg_bank[846] ,
         \iRF_stage/reg_bank/reg_bank[847] ,
         \iRF_stage/reg_bank/reg_bank[848] ,
         \iRF_stage/reg_bank/reg_bank[849] ,
         \iRF_stage/reg_bank/reg_bank[850] ,
         \iRF_stage/reg_bank/reg_bank[851] ,
         \iRF_stage/reg_bank/reg_bank[852] ,
         \iRF_stage/reg_bank/reg_bank[853] ,
         \iRF_stage/reg_bank/reg_bank[854] ,
         \iRF_stage/reg_bank/reg_bank[855] ,
         \iRF_stage/reg_bank/reg_bank[856] ,
         \iRF_stage/reg_bank/reg_bank[857] ,
         \iRF_stage/reg_bank/reg_bank[858] ,
         \iRF_stage/reg_bank/reg_bank[859] ,
         \iRF_stage/reg_bank/reg_bank[860] ,
         \iRF_stage/reg_bank/reg_bank[861] ,
         \iRF_stage/reg_bank/reg_bank[862] ,
         \iRF_stage/reg_bank/reg_bank[863] ,
         \iRF_stage/reg_bank/reg_bank[864] ,
         \iRF_stage/reg_bank/reg_bank[865] ,
         \iRF_stage/reg_bank/reg_bank[866] ,
         \iRF_stage/reg_bank/reg_bank[867] ,
         \iRF_stage/reg_bank/reg_bank[868] ,
         \iRF_stage/reg_bank/reg_bank[869] ,
         \iRF_stage/reg_bank/reg_bank[870] ,
         \iRF_stage/reg_bank/reg_bank[871] ,
         \iRF_stage/reg_bank/reg_bank[872] ,
         \iRF_stage/reg_bank/reg_bank[873] ,
         \iRF_stage/reg_bank/reg_bank[874] ,
         \iRF_stage/reg_bank/reg_bank[875] ,
         \iRF_stage/reg_bank/reg_bank[876] ,
         \iRF_stage/reg_bank/reg_bank[877] ,
         \iRF_stage/reg_bank/reg_bank[878] ,
         \iRF_stage/reg_bank/reg_bank[879] ,
         \iRF_stage/reg_bank/reg_bank[880] ,
         \iRF_stage/reg_bank/reg_bank[881] ,
         \iRF_stage/reg_bank/reg_bank[882] ,
         \iRF_stage/reg_bank/reg_bank[883] ,
         \iRF_stage/reg_bank/reg_bank[884] ,
         \iRF_stage/reg_bank/reg_bank[885] ,
         \iRF_stage/reg_bank/reg_bank[886] ,
         \iRF_stage/reg_bank/reg_bank[887] ,
         \iRF_stage/reg_bank/reg_bank[888] ,
         \iRF_stage/reg_bank/reg_bank[889] ,
         \iRF_stage/reg_bank/reg_bank[890] ,
         \iRF_stage/reg_bank/reg_bank[891] ,
         \iRF_stage/reg_bank/reg_bank[892] ,
         \iRF_stage/reg_bank/reg_bank[893] ,
         \iRF_stage/reg_bank/reg_bank[894] ,
         \iRF_stage/reg_bank/reg_bank[895] ,
         \iRF_stage/reg_bank/reg_bank[896] ,
         \iRF_stage/reg_bank/reg_bank[897] ,
         \iRF_stage/reg_bank/reg_bank[898] ,
         \iRF_stage/reg_bank/reg_bank[899] ,
         \iRF_stage/reg_bank/reg_bank[900] ,
         \iRF_stage/reg_bank/reg_bank[901] ,
         \iRF_stage/reg_bank/reg_bank[902] ,
         \iRF_stage/reg_bank/reg_bank[903] ,
         \iRF_stage/reg_bank/reg_bank[904] ,
         \iRF_stage/reg_bank/reg_bank[905] ,
         \iRF_stage/reg_bank/reg_bank[906] ,
         \iRF_stage/reg_bank/reg_bank[907] ,
         \iRF_stage/reg_bank/reg_bank[908] ,
         \iRF_stage/reg_bank/reg_bank[909] ,
         \iRF_stage/reg_bank/reg_bank[910] ,
         \iRF_stage/reg_bank/reg_bank[911] ,
         \iRF_stage/reg_bank/reg_bank[912] ,
         \iRF_stage/reg_bank/reg_bank[913] ,
         \iRF_stage/reg_bank/reg_bank[914] ,
         \iRF_stage/reg_bank/reg_bank[915] ,
         \iRF_stage/reg_bank/reg_bank[916] ,
         \iRF_stage/reg_bank/reg_bank[917] ,
         \iRF_stage/reg_bank/reg_bank[918] ,
         \iRF_stage/reg_bank/reg_bank[919] ,
         \iRF_stage/reg_bank/reg_bank[920] ,
         \iRF_stage/reg_bank/reg_bank[921] ,
         \iRF_stage/reg_bank/reg_bank[922] ,
         \iRF_stage/reg_bank/reg_bank[923] ,
         \iRF_stage/reg_bank/reg_bank[924] ,
         \iRF_stage/reg_bank/reg_bank[925] ,
         \iRF_stage/reg_bank/reg_bank[926] ,
         \iRF_stage/reg_bank/reg_bank[927] ,
         \iRF_stage/reg_bank/reg_bank[928] ,
         \iRF_stage/reg_bank/reg_bank[929] ,
         \iRF_stage/reg_bank/reg_bank[930] ,
         \iRF_stage/reg_bank/reg_bank[931] ,
         \iRF_stage/reg_bank/reg_bank[932] ,
         \iRF_stage/reg_bank/reg_bank[933] ,
         \iRF_stage/reg_bank/reg_bank[934] ,
         \iRF_stage/reg_bank/reg_bank[935] ,
         \iRF_stage/reg_bank/reg_bank[936] ,
         \iRF_stage/reg_bank/reg_bank[937] ,
         \iRF_stage/reg_bank/reg_bank[938] ,
         \iRF_stage/reg_bank/reg_bank[939] ,
         \iRF_stage/reg_bank/reg_bank[940] ,
         \iRF_stage/reg_bank/reg_bank[941] ,
         \iRF_stage/reg_bank/reg_bank[942] ,
         \iRF_stage/reg_bank/reg_bank[943] ,
         \iRF_stage/reg_bank/reg_bank[944] ,
         \iRF_stage/reg_bank/reg_bank[945] ,
         \iRF_stage/reg_bank/reg_bank[946] ,
         \iRF_stage/reg_bank/reg_bank[947] ,
         \iRF_stage/reg_bank/reg_bank[948] ,
         \iRF_stage/reg_bank/reg_bank[949] ,
         \iRF_stage/reg_bank/reg_bank[950] ,
         \iRF_stage/reg_bank/reg_bank[951] ,
         \iRF_stage/reg_bank/reg_bank[952] ,
         \iRF_stage/reg_bank/reg_bank[953] ,
         \iRF_stage/reg_bank/reg_bank[954] ,
         \iRF_stage/reg_bank/reg_bank[955] ,
         \iRF_stage/reg_bank/reg_bank[956] ,
         \iRF_stage/reg_bank/reg_bank[957] ,
         \iRF_stage/reg_bank/reg_bank[958] ,
         \iRF_stage/reg_bank/reg_bank[959] ,
         \iRF_stage/reg_bank/reg_bank[960] ,
         \iRF_stage/reg_bank/reg_bank[961] ,
         \iRF_stage/reg_bank/reg_bank[962] ,
         \iRF_stage/reg_bank/reg_bank[963] ,
         \iRF_stage/reg_bank/reg_bank[964] ,
         \iRF_stage/reg_bank/reg_bank[965] ,
         \iRF_stage/reg_bank/reg_bank[966] ,
         \iRF_stage/reg_bank/reg_bank[967] ,
         \iRF_stage/reg_bank/reg_bank[968] ,
         \iRF_stage/reg_bank/reg_bank[969] ,
         \iRF_stage/reg_bank/reg_bank[970] ,
         \iRF_stage/reg_bank/reg_bank[971] ,
         \iRF_stage/reg_bank/reg_bank[972] ,
         \iRF_stage/reg_bank/reg_bank[973] ,
         \iRF_stage/reg_bank/reg_bank[974] ,
         \iRF_stage/reg_bank/reg_bank[975] ,
         \iRF_stage/reg_bank/reg_bank[976] ,
         \iRF_stage/reg_bank/reg_bank[977] ,
         \iRF_stage/reg_bank/reg_bank[978] ,
         \iRF_stage/reg_bank/reg_bank[979] ,
         \iRF_stage/reg_bank/reg_bank[980] ,
         \iRF_stage/reg_bank/reg_bank[981] ,
         \iRF_stage/reg_bank/reg_bank[982] ,
         \iRF_stage/reg_bank/reg_bank[983] ,
         \iRF_stage/reg_bank/reg_bank[984] ,
         \iRF_stage/reg_bank/reg_bank[985] ,
         \iRF_stage/reg_bank/reg_bank[986] ,
         \iRF_stage/reg_bank/reg_bank[987] ,
         \iRF_stage/reg_bank/reg_bank[988] ,
         \iRF_stage/reg_bank/reg_bank[989] ,
         \iRF_stage/reg_bank/reg_bank[990] ,
         \iRF_stage/reg_bank/reg_bank[991] ,
         \iRF_stage/reg_bank/reg_bank[992] ,
         \iRF_stage/reg_bank/reg_bank[993] ,
         \iRF_stage/reg_bank/reg_bank[994] ,
         \iRF_stage/reg_bank/reg_bank[995] ,
         \iRF_stage/reg_bank/reg_bank[996] ,
         \iRF_stage/reg_bank/reg_bank[997] ,
         \iRF_stage/reg_bank/reg_bank[998] ,
         \iRF_stage/reg_bank/reg_bank[999] ,
         \iRF_stage/reg_bank/reg_bank[1000] ,
         \iRF_stage/reg_bank/reg_bank[1001] ,
         \iRF_stage/reg_bank/reg_bank[1002] ,
         \iRF_stage/reg_bank/reg_bank[1003] ,
         \iRF_stage/reg_bank/reg_bank[1004] ,
         \iRF_stage/reg_bank/reg_bank[1005] ,
         \iRF_stage/reg_bank/reg_bank[1006] ,
         \iRF_stage/reg_bank/reg_bank[1007] ,
         \iRF_stage/reg_bank/reg_bank[1008] ,
         \iRF_stage/reg_bank/reg_bank[1009] ,
         \iRF_stage/reg_bank/reg_bank[1010] ,
         \iRF_stage/reg_bank/reg_bank[1011] ,
         \iRF_stage/reg_bank/reg_bank[1012] ,
         \iRF_stage/reg_bank/reg_bank[1013] ,
         \iRF_stage/reg_bank/reg_bank[1014] ,
         \iRF_stage/reg_bank/reg_bank[1015] ,
         \iRF_stage/reg_bank/reg_bank[1016] ,
         \iRF_stage/reg_bank/reg_bank[1017] ,
         \iRF_stage/reg_bank/reg_bank[1018] ,
         \iRF_stage/reg_bank/reg_bank[1019] ,
         \iRF_stage/reg_bank/reg_bank[1020] ,
         \iRF_stage/reg_bank/reg_bank[1021] ,
         \iRF_stage/reg_bank/reg_bank[1022] ,
         \iRF_stage/reg_bank/reg_bank[1023] , \iRF_stage/reg_bank/r_wren ,
         \iRF_stage/reg_bank/r_wraddress[0] ,
         \iRF_stage/reg_bank/r_wraddress[1] ,
         \iRF_stage/reg_bank/r_wraddress[2] ,
         \iRF_stage/reg_bank/r_wraddress[3] ,
         \iRF_stage/reg_bank/r_wraddress[4] , \iRF_stage/reg_bank/N21 ,
         \iRF_stage/reg_bank/N20 , \iRF_stage/reg_bank/N19 ,
         \iRF_stage/reg_bank/N18 , \iRF_stage/reg_bank/N17 ,
         \iRF_stage/reg_bank/N16 , \iRF_stage/reg_bank/N15 ,
         \iRF_stage/reg_bank/N14 , \iRF_stage/reg_bank/N13 ,
         \iRF_stage/reg_bank/N12 , \decoder_pipe/pipereg/BUS4987[0] ,
         \decoder_pipe/pipereg/BUS7299[0] , \decoder_pipe/pipereg/BUS7822[0] ,
         \decoder_pipe/pipereg/BUS5682[0] , \decoder_pipe/pipereg/BUS5790[0] ,
         \decoder_pipe/pipereg/BUS5008[1] , \decoder_pipe/pipereg/BUS5008[0] ,
         \decoder_pipe/pipereg/BUS5674[4] , \decoder_pipe/pipereg/BUS5674[3] ,
         \decoder_pipe/pipereg/BUS5674[2] , \decoder_pipe/pipereg/BUS5674[1] ,
         \decoder_pipe/pipereg/BUS5674[0] , \decoder_pipe/pipereg/BUS5666[3] ,
         \decoder_pipe/pipereg/BUS5666[2] , \decoder_pipe/pipereg/BUS5666[1] ,
         \decoder_pipe/pipereg/BUS5666[0] , \decoder_pipe/pipereg/BUS5690[0] ,
         \decoder_pipe/pipereg/NET7643 , \decoder_pipe/pipereg/BUS5639[0] ,
         \decoder_pipe/pipereg/BUS5651[0] , \decoder_pipe/pipereg/BUS5483[1] ,
         \decoder_pipe/pipereg/BUS5483[0] ,
         \iexec_stage/MIPS_alu/mips_shifter/n601 ,
         \iexec_stage/MIPS_alu/mips_shifter/n600 ,
         \iexec_stage/MIPS_alu/mips_shifter/n598 ,
         \iexec_stage/MIPS_alu/mips_shifter/n597 ,
         \iexec_stage/MIPS_alu/mips_shifter/n596 ,
         \iexec_stage/MIPS_alu/mips_shifter/n595 ,
         \iexec_stage/MIPS_alu/mips_shifter/n593 ,
         \iexec_stage/MIPS_alu/mips_shifter/n592 ,
         \iexec_stage/MIPS_alu/mips_shifter/n590 ,
         \iexec_stage/MIPS_alu/mips_shifter/n589 ,
         \iexec_stage/MIPS_alu/mips_shifter/n588 ,
         \iexec_stage/MIPS_alu/mips_shifter/n586 ,
         \iexec_stage/MIPS_alu/mips_shifter/n585 ,
         \iexec_stage/MIPS_alu/mips_shifter/n584 ,
         \iexec_stage/MIPS_alu/mips_shifter/n582 ,
         \iexec_stage/MIPS_alu/mips_shifter/n581 ,
         \iexec_stage/MIPS_alu/mips_shifter/n580 ,
         \iexec_stage/MIPS_alu/mips_shifter/n578 ,
         \iexec_stage/MIPS_alu/mips_shifter/n577 ,
         \iexec_stage/MIPS_alu/mips_shifter/n576 ,
         \iexec_stage/MIPS_alu/mips_shifter/n574 ,
         \iexec_stage/MIPS_alu/mips_shifter/n573 ,
         \iexec_stage/MIPS_alu/mips_shifter/n572 ,
         \iexec_stage/MIPS_alu/mips_shifter/n570 ,
         \iexec_stage/MIPS_alu/mips_shifter/n569 ,
         \iexec_stage/MIPS_alu/mips_shifter/n568 ,
         \iexec_stage/MIPS_alu/mips_shifter/n565 ,
         \iexec_stage/MIPS_alu/mips_shifter/n564 ,
         \iexec_stage/MIPS_alu/mips_shifter/n562 ,
         \iexec_stage/MIPS_alu/mips_shifter/n560 ,
         \iexec_stage/MIPS_alu/mips_shifter/n559 ,
         \iexec_stage/MIPS_alu/mips_shifter/n558 ,
         \iexec_stage/MIPS_alu/mips_shifter/n557 ,
         \iexec_stage/MIPS_alu/mips_shifter/n556 ,
         \iexec_stage/MIPS_alu/mips_shifter/n555 ,
         \iexec_stage/MIPS_alu/mips_shifter/n553 ,
         \iexec_stage/MIPS_alu/mips_shifter/n552 ,
         \iexec_stage/MIPS_alu/mips_shifter/n551 ,
         \iexec_stage/MIPS_alu/mips_shifter/n550 ,
         \iexec_stage/MIPS_alu/mips_shifter/n549 ,
         \iexec_stage/MIPS_alu/mips_shifter/n548 ,
         \iexec_stage/MIPS_alu/mips_shifter/n546 ,
         \iexec_stage/MIPS_alu/mips_shifter/n545 ,
         \iexec_stage/MIPS_alu/mips_shifter/n544 ,
         \iexec_stage/MIPS_alu/mips_shifter/n543 ,
         \iexec_stage/MIPS_alu/mips_shifter/n542 ,
         \iexec_stage/MIPS_alu/mips_shifter/n541 ,
         \iexec_stage/MIPS_alu/mips_shifter/n540 ,
         \iexec_stage/MIPS_alu/mips_shifter/n539 ,
         \iexec_stage/MIPS_alu/mips_shifter/n538 ,
         \iexec_stage/MIPS_alu/mips_shifter/n537 ,
         \iexec_stage/MIPS_alu/mips_shifter/n536 ,
         \iexec_stage/MIPS_alu/mips_shifter/n535 ,
         \iexec_stage/MIPS_alu/mips_shifter/n534 ,
         \iexec_stage/MIPS_alu/mips_shifter/n530 ,
         \iexec_stage/MIPS_alu/mips_shifter/n528 ,
         \iexec_stage/MIPS_alu/mips_shifter/n526 ,
         \iexec_stage/MIPS_alu/mips_shifter/n524 ,
         \iexec_stage/MIPS_alu/mips_shifter/n522 ,
         \iexec_stage/MIPS_alu/mips_shifter/n520 ,
         \iexec_stage/MIPS_alu/mips_shifter/n519 ,
         \iexec_stage/MIPS_alu/mips_shifter/n518 ,
         \iexec_stage/MIPS_alu/mips_shifter/n516 ,
         \iexec_stage/MIPS_alu/mips_shifter/n515 ,
         \iexec_stage/MIPS_alu/mips_shifter/n514 ,
         \iexec_stage/MIPS_alu/mips_shifter/n512 ,
         \iexec_stage/MIPS_alu/mips_shifter/n511 ,
         \iexec_stage/MIPS_alu/mips_shifter/n510 ,
         \iexec_stage/MIPS_alu/mips_shifter/n509 ,
         \iexec_stage/MIPS_alu/mips_shifter/n508 ,
         \iexec_stage/MIPS_alu/mips_shifter/n507 ,
         \iexec_stage/MIPS_alu/mips_shifter/n505 ,
         \iexec_stage/MIPS_alu/mips_shifter/n504 ,
         \iexec_stage/MIPS_alu/mips_shifter/n503 ,
         \iexec_stage/MIPS_alu/mips_shifter/n501 ,
         \iexec_stage/MIPS_alu/mips_shifter/n500 ,
         \iexec_stage/MIPS_alu/mips_shifter/n499 ,
         \iexec_stage/MIPS_alu/mips_shifter/n497 ,
         \iexec_stage/MIPS_alu/mips_shifter/n496 ,
         \iexec_stage/MIPS_alu/mips_shifter/n495 ,
         \iexec_stage/MIPS_alu/mips_shifter/n493 ,
         \iexec_stage/MIPS_alu/mips_shifter/n492 ,
         \iexec_stage/MIPS_alu/mips_shifter/n491 ,
         \iexec_stage/MIPS_alu/mips_shifter/n489 ,
         \iexec_stage/MIPS_alu/mips_shifter/n488 ,
         \iexec_stage/MIPS_alu/mips_shifter/n487 ,
         \iexec_stage/MIPS_alu/mips_shifter/n485 ,
         \iexec_stage/MIPS_alu/mips_shifter/n484 ,
         \iexec_stage/MIPS_alu/mips_shifter/n483 ,
         \iexec_stage/MIPS_alu/mips_shifter/n481 ,
         \iexec_stage/MIPS_alu/mips_shifter/n480 ,
         \iexec_stage/MIPS_alu/mips_shifter/n479 ,
         \iexec_stage/MIPS_alu/mips_shifter/n478 ,
         \iexec_stage/MIPS_alu/mips_shifter/n477 ,
         \iexec_stage/MIPS_alu/mips_shifter/n476 ,
         \iexec_stage/MIPS_alu/mips_shifter/n475 ,
         \iexec_stage/MIPS_alu/mips_shifter/n473 ,
         \iexec_stage/MIPS_alu/mips_shifter/n472 ,
         \iexec_stage/MIPS_alu/mips_shifter/n471 ,
         \iexec_stage/MIPS_alu/mips_shifter/n470 ,
         \iexec_stage/MIPS_alu/mips_shifter/n468 ,
         \iexec_stage/MIPS_alu/mips_shifter/n467 ,
         \iexec_stage/MIPS_alu/mips_shifter/n466 ,
         \iexec_stage/MIPS_alu/mips_shifter/n465 ,
         \iexec_stage/MIPS_alu/mips_shifter/n463 ,
         \iexec_stage/MIPS_alu/mips_shifter/n462 ,
         \iexec_stage/MIPS_alu/mips_shifter/n461 ,
         \iexec_stage/MIPS_alu/mips_shifter/n460 ,
         \iexec_stage/MIPS_alu/mips_shifter/n458 ,
         \iexec_stage/MIPS_alu/mips_shifter/n457 ,
         \iexec_stage/MIPS_alu/mips_shifter/n456 ,
         \iexec_stage/MIPS_alu/mips_shifter/n455 ,
         \iexec_stage/MIPS_alu/mips_shifter/n453 ,
         \iexec_stage/MIPS_alu/mips_shifter/n452 ,
         \iexec_stage/MIPS_alu/mips_shifter/n451 ,
         \iexec_stage/MIPS_alu/mips_shifter/n450 ,
         \iexec_stage/MIPS_alu/mips_shifter/n449 ,
         \iexec_stage/MIPS_alu/mips_shifter/n447 ,
         \iexec_stage/MIPS_alu/mips_shifter/n446 ,
         \iexec_stage/MIPS_alu/mips_shifter/n445 ,
         \iexec_stage/MIPS_alu/mips_shifter/n444 ,
         \iexec_stage/MIPS_alu/mips_shifter/n443 ,
         \iexec_stage/MIPS_alu/mips_shifter/n442 ,
         \iexec_stage/MIPS_alu/mips_shifter/n441 ,
         \iexec_stage/MIPS_alu/mips_shifter/n440 ,
         \iexec_stage/MIPS_alu/mips_shifter/n439 ,
         \iexec_stage/MIPS_alu/mips_shifter/n438 ,
         \iexec_stage/MIPS_alu/mips_shifter/n437 ,
         \iexec_stage/MIPS_alu/mips_shifter/n436 ,
         \iexec_stage/MIPS_alu/mips_shifter/n435 ,
         \iexec_stage/MIPS_alu/mips_shifter/n434 ,
         \iexec_stage/MIPS_alu/mips_shifter/n431 ,
         \iexec_stage/MIPS_alu/mips_shifter/n430 ,
         \iexec_stage/MIPS_alu/mips_shifter/n429 ,
         \iexec_stage/MIPS_alu/mips_shifter/n427 ,
         \iexec_stage/MIPS_alu/mips_shifter/n426 ,
         \iexec_stage/MIPS_alu/mips_shifter/n425 ,
         \iexec_stage/MIPS_alu/mips_shifter/n422 ,
         \iexec_stage/MIPS_alu/mips_shifter/n419 ,
         \iexec_stage/MIPS_alu/mips_shifter/n418 ,
         \iexec_stage/MIPS_alu/mips_shifter/n417 ,
         \iexec_stage/MIPS_alu/mips_shifter/n416 ,
         \iexec_stage/MIPS_alu/mips_shifter/n415 ,
         \iexec_stage/MIPS_alu/mips_shifter/n414 ,
         \iexec_stage/MIPS_alu/mips_shifter/n413 ,
         \iexec_stage/MIPS_alu/mips_shifter/n412 ,
         \iexec_stage/MIPS_alu/mips_shifter/n411 ,
         \iexec_stage/MIPS_alu/mips_shifter/n410 ,
         \iexec_stage/MIPS_alu/mips_shifter/n409 ,
         \iexec_stage/MIPS_alu/mips_shifter/n408 ,
         \iexec_stage/MIPS_alu/mips_shifter/n407 ,
         \iexec_stage/MIPS_alu/mips_shifter/n405 ,
         \iexec_stage/MIPS_alu/mips_shifter/n404 ,
         \iexec_stage/MIPS_alu/mips_shifter/n403 ,
         \iexec_stage/MIPS_alu/mips_shifter/n402 ,
         \iexec_stage/MIPS_alu/mips_shifter/n401 ,
         \iexec_stage/MIPS_alu/mips_shifter/n400 ,
         \iexec_stage/MIPS_alu/mips_shifter/n399 ,
         \iexec_stage/MIPS_alu/mips_shifter/n398 ,
         \iexec_stage/MIPS_alu/mips_shifter/n397 ,
         \iexec_stage/MIPS_alu/mips_shifter/n396 ,
         \iexec_stage/MIPS_alu/mips_shifter/n395 ,
         \iexec_stage/MIPS_alu/mips_shifter/n394 ,
         \iexec_stage/MIPS_alu/mips_shifter/n393 ,
         \iexec_stage/MIPS_alu/mips_shifter/n392 ,
         \iexec_stage/MIPS_alu/mips_shifter/n391 ,
         \iexec_stage/MIPS_alu/mips_shifter/n390 ,
         \iexec_stage/MIPS_alu/mips_shifter/n389 ,
         \iexec_stage/MIPS_alu/mips_shifter/n388 ,
         \iexec_stage/MIPS_alu/mips_shifter/n387 ,
         \iexec_stage/MIPS_alu/mips_shifter/n386 ,
         \iexec_stage/MIPS_alu/mips_shifter/n385 ,
         \iexec_stage/MIPS_alu/mips_shifter/n384 ,
         \iexec_stage/MIPS_alu/mips_shifter/n383 ,
         \iexec_stage/MIPS_alu/mips_shifter/n382 ,
         \iexec_stage/MIPS_alu/mips_shifter/n381 ,
         \iexec_stage/MIPS_alu/mips_shifter/n380 ,
         \iexec_stage/MIPS_alu/mips_shifter/n378 ,
         \iexec_stage/MIPS_alu/mips_shifter/n377 ,
         \iexec_stage/MIPS_alu/mips_shifter/n376 ,
         \iexec_stage/MIPS_alu/mips_shifter/n375 ,
         \iexec_stage/MIPS_alu/mips_shifter/n374 ,
         \iexec_stage/MIPS_alu/mips_shifter/n373 ,
         \iexec_stage/MIPS_alu/mips_shifter/n372 ,
         \iexec_stage/MIPS_alu/mips_shifter/n370 ,
         \iexec_stage/MIPS_alu/mips_shifter/n369 ,
         \iexec_stage/MIPS_alu/mips_shifter/n368 ,
         \iexec_stage/MIPS_alu/mips_shifter/n367 ,
         \iexec_stage/MIPS_alu/mips_shifter/n366 ,
         \iexec_stage/MIPS_alu/mips_shifter/n365 ,
         \iexec_stage/MIPS_alu/mips_shifter/n364 ,
         \iexec_stage/MIPS_alu/mips_shifter/n363 ,
         \iexec_stage/MIPS_alu/mips_shifter/n362 ,
         \iexec_stage/MIPS_alu/mips_shifter/n361 ,
         \iexec_stage/MIPS_alu/mips_shifter/n360 ,
         \iexec_stage/MIPS_alu/mips_shifter/n359 ,
         \iexec_stage/MIPS_alu/mips_shifter/N256 ,
         \iexec_stage/MIPS_alu/mips_shifter/N255 ,
         \iexec_stage/MIPS_alu/mips_shifter/N254 ,
         \iexec_stage/MIPS_alu/mips_shifter/N253 ,
         \iexec_stage/MIPS_alu/mips_shifter/N252 ,
         \iexec_stage/MIPS_alu/mips_shifter/N251 ,
         \iexec_stage/MIPS_alu/mips_shifter/N250 ,
         \iexec_stage/MIPS_alu/mips_shifter/N249 ,
         \iexec_stage/MIPS_alu/mips_shifter/N248 ,
         \iexec_stage/MIPS_alu/mips_shifter/N247 ,
         \iexec_stage/MIPS_alu/mips_shifter/N246 ,
         \iexec_stage/MIPS_alu/mips_shifter/N245 ,
         \iexec_stage/MIPS_alu/mips_shifter/N244 ,
         \iexec_stage/MIPS_alu/mips_shifter/N243 ,
         \iexec_stage/MIPS_alu/mips_shifter/N242 ,
         \iexec_stage/MIPS_alu/mips_shifter/N224 ,
         \iexec_stage/MIPS_alu/mips_shifter/N223 ,
         \iexec_stage/MIPS_alu/mips_shifter/N222 ,
         \iexec_stage/MIPS_alu/mips_shifter/N221 ,
         \iexec_stage/MIPS_alu/mips_shifter/N220 ,
         \iexec_stage/MIPS_alu/mips_shifter/N219 ,
         \iexec_stage/MIPS_alu/mips_shifter/N218 ,
         \iexec_stage/MIPS_alu/mips_shifter/N217 ,
         \iexec_stage/MIPS_alu/mips_shifter/N216 ,
         \iexec_stage/MIPS_alu/mips_shifter/N215 ,
         \iexec_stage/MIPS_alu/mips_shifter/N214 ,
         \iexec_stage/MIPS_alu/mips_shifter/N213 ,
         \iexec_stage/MIPS_alu/mips_shifter/N212 ,
         \iexec_stage/MIPS_alu/mips_shifter/N211 ,
         \iexec_stage/MIPS_alu/mips_shifter/N210 ,
         \iexec_stage/MIPS_alu/mips_shifter/N208 ,
         \iexec_stage/MIPS_alu/mips_shifter/N207 ,
         \iexec_stage/MIPS_alu/mips_shifter/N206 ,
         \iexec_stage/MIPS_alu/mips_shifter/N205 ,
         \iexec_stage/MIPS_alu/mips_shifter/N204 ,
         \iexec_stage/MIPS_alu/mips_shifter/N203 ,
         \iexec_stage/MIPS_alu/mips_shifter/N202 ,
         \iexec_stage/MIPS_alu/mips_shifter/N201 ,
         \iexec_stage/MIPS_alu/mips_shifter/N200 ,
         \iexec_stage/MIPS_alu/mips_shifter/N199 ,
         \iexec_stage/MIPS_alu/mips_shifter/N198 ,
         \iexec_stage/MIPS_alu/mips_shifter/N197 ,
         \iexec_stage/MIPS_alu/mips_shifter/N196 ,
         \iexec_stage/MIPS_alu/mips_shifter/N195 ,
         \iexec_stage/MIPS_alu/mips_shifter/N194 ,
         \iexec_stage/MIPS_alu/mips_shifter/N193 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_32 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_30 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_29 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_28 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_27 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_26 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_25 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_24 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_23 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_22 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_21 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_20 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_19 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_18 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_17 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_16 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_15 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_14 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_13 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_12 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_11 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_10 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_9 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_8 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_7 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_6 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_5 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_4 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_3 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_2 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_1 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_0 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_32 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_30 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_29 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_28 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_27 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_26 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_25 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_24 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_23 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_22 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_21 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_20 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_19 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_18 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_17 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_16 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_15 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_14 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_13 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_12 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_11 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_10 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_9 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_8 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_7 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_6 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_5 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_4 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_3 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_2 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_1 ,
         \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_0 ,
         \iexec_stage/MIPS_alu/mips_alu/N370 ,
         \iexec_stage/MIPS_alu/mips_alu/N207 ,
         \iexec_stage/MIPS_alu/mips_alu/N206 ,
         \iexec_stage/MIPS_alu/mips_alu/N205 ,
         \iexec_stage/MIPS_alu/mips_alu/N204 ,
         \iexec_stage/MIPS_alu/mips_alu/N203 ,
         \iexec_stage/MIPS_alu/mips_alu/N202 ,
         \iexec_stage/MIPS_alu/mips_alu/N201 ,
         \iexec_stage/MIPS_alu/mips_alu/N200 ,
         \iexec_stage/MIPS_alu/mips_alu/N199 ,
         \iexec_stage/MIPS_alu/mips_alu/N198 ,
         \iexec_stage/MIPS_alu/mips_alu/N197 ,
         \iexec_stage/MIPS_alu/mips_alu/N196 ,
         \iexec_stage/MIPS_alu/mips_alu/N195 ,
         \iexec_stage/MIPS_alu/mips_alu/N194 ,
         \iexec_stage/MIPS_alu/mips_alu/N193 ,
         \iexec_stage/MIPS_alu/mips_alu/N192 ,
         \iexec_stage/MIPS_alu/mips_alu/N191 ,
         \iexec_stage/MIPS_alu/mips_alu/N190 ,
         \iexec_stage/MIPS_alu/mips_alu/N189 ,
         \iexec_stage/MIPS_alu/mips_alu/N188 ,
         \iexec_stage/MIPS_alu/mips_alu/N187 ,
         \iexec_stage/MIPS_alu/mips_alu/N186 ,
         \iexec_stage/MIPS_alu/mips_alu/N185 ,
         \iexec_stage/MIPS_alu/mips_alu/N184 ,
         \iexec_stage/MIPS_alu/mips_alu/N183 ,
         \iexec_stage/MIPS_alu/mips_alu/N182 ,
         \iexec_stage/MIPS_alu/mips_alu/N181 ,
         \iexec_stage/MIPS_alu/mips_alu/N180 ,
         \iexec_stage/MIPS_alu/mips_alu/N179 ,
         \iexec_stage/MIPS_alu/mips_alu/N178 ,
         \iexec_stage/MIPS_alu/mips_alu/N177 ,
         \iexec_stage/MIPS_alu/mips_alu/N176 ,
         \iexec_stage/MIPS_alu/mips_alu/N143 ,
         \iexec_stage/MIPS_alu/mips_alu/N142 ,
         \iexec_stage/MIPS_alu/mips_alu/N141 ,
         \iexec_stage/MIPS_alu/mips_alu/N140 ,
         \iexec_stage/MIPS_alu/mips_alu/N139 ,
         \iexec_stage/MIPS_alu/mips_alu/N138 ,
         \iexec_stage/MIPS_alu/mips_alu/N137 ,
         \iexec_stage/MIPS_alu/mips_alu/N136 ,
         \iexec_stage/MIPS_alu/mips_alu/N135 ,
         \iexec_stage/MIPS_alu/mips_alu/N134 ,
         \iexec_stage/MIPS_alu/mips_alu/N133 ,
         \iexec_stage/MIPS_alu/mips_alu/N132 ,
         \iexec_stage/MIPS_alu/mips_alu/N131 ,
         \iexec_stage/MIPS_alu/mips_alu/N130 ,
         \iexec_stage/MIPS_alu/mips_alu/N129 ,
         \iexec_stage/MIPS_alu/mips_alu/N128 ,
         \iexec_stage/MIPS_alu/mips_alu/N127 ,
         \iexec_stage/MIPS_alu/mips_alu/N126 ,
         \iexec_stage/MIPS_alu/mips_alu/N125 ,
         \iexec_stage/MIPS_alu/mips_alu/N124 ,
         \iexec_stage/MIPS_alu/mips_alu/N123 ,
         \iexec_stage/MIPS_alu/mips_alu/N122 ,
         \iexec_stage/MIPS_alu/mips_alu/N121 ,
         \iexec_stage/MIPS_alu/mips_alu/N120 ,
         \iexec_stage/MIPS_alu/mips_alu/N119 ,
         \iexec_stage/MIPS_alu/mips_alu/N118 ,
         \iexec_stage/MIPS_alu/mips_alu/N117 ,
         \iexec_stage/MIPS_alu/mips_alu/N116 ,
         \iexec_stage/MIPS_alu/mips_alu/N115 ,
         \iexec_stage/MIPS_alu/mips_alu/N114 ,
         \iexec_stage/MIPS_alu/mips_alu/N113 ,
         \iexec_stage/MIPS_alu/mips_alu/N112 , \decoder_pipe/pipereg/U10/n4 ,
         \decoder_pipe/pipereg/U11/n4 , \decoder_pipe/pipereg/U6/n4 ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[31] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[30] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[29] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[28] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[27] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[26] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[25] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[24] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[23] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[22] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[21] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[20] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[19] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[18] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[17] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[16] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[15] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[14] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[13] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[12] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[11] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[10] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[9] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[8] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[7] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[6] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[5] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[4] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[3] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[2] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[1] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[0] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[1] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[2] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[3] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[4] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[5] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[6] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[7] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[8] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[9] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[10] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[11] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[12] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[13] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[14] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[15] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[16] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[17] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[18] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[19] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[20] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[21] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[22] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[23] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[24] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[25] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[26] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[27] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[28] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[29] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[30] ,
         \iexec_stage/MIPS_alu/mips_alu/r92/carry[31] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[32] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[31] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[30] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[29] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[28] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[27] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[26] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[25] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[24] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[23] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[22] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[21] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[20] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[19] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[18] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[17] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[16] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[15] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[14] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[13] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[12] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[11] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[10] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[9] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[8] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[7] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[6] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[5] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[4] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[3] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[2] ,
         \iexec_stage/MIPS_alu/mips_alu/r86/carry[1] ,
         \iexec_stage/add4/add_39/carry[31] ,
         \iexec_stage/add4/add_39/carry[30] ,
         \iexec_stage/add4/add_39/carry[29] ,
         \iexec_stage/add4/add_39/carry[28] ,
         \iexec_stage/add4/add_39/carry[27] ,
         \iexec_stage/add4/add_39/carry[26] ,
         \iexec_stage/add4/add_39/carry[25] ,
         \iexec_stage/add4/add_39/carry[24] ,
         \iexec_stage/add4/add_39/carry[23] ,
         \iexec_stage/add4/add_39/carry[22] ,
         \iexec_stage/add4/add_39/carry[21] ,
         \iexec_stage/add4/add_39/carry[20] ,
         \iexec_stage/add4/add_39/carry[19] ,
         \iexec_stage/add4/add_39/carry[18] ,
         \iexec_stage/add4/add_39/carry[17] ,
         \iexec_stage/add4/add_39/carry[16] ,
         \iexec_stage/add4/add_39/carry[15] ,
         \iexec_stage/add4/add_39/carry[14] ,
         \iexec_stage/add4/add_39/carry[13] ,
         \iexec_stage/add4/add_39/carry[12] ,
         \iexec_stage/add4/add_39/carry[11] ,
         \iexec_stage/add4/add_39/carry[10] ,
         \iexec_stage/add4/add_39/carry[9] ,
         \iexec_stage/add4/add_39/carry[8] ,
         \iexec_stage/add4/add_39/carry[7] ,
         \iexec_stage/add4/add_39/carry[6] ,
         \iexec_stage/add4/add_39/carry[5] ,
         \iexec_stage/add4/add_39/carry[4] ,
         \iRF_stage/i_pc_gen/r62/carry[31] ,
         \iRF_stage/i_pc_gen/r62/carry[30] ,
         \iRF_stage/i_pc_gen/r62/carry[29] ,
         \iRF_stage/i_pc_gen/r62/carry[28] ,
         \iRF_stage/i_pc_gen/r62/carry[27] ,
         \iRF_stage/i_pc_gen/r62/carry[26] ,
         \iRF_stage/i_pc_gen/r62/carry[25] ,
         \iRF_stage/i_pc_gen/r62/carry[24] ,
         \iRF_stage/i_pc_gen/r62/carry[23] ,
         \iRF_stage/i_pc_gen/r62/carry[22] ,
         \iRF_stage/i_pc_gen/r62/carry[21] ,
         \iRF_stage/i_pc_gen/r62/carry[20] ,
         \iRF_stage/i_pc_gen/r62/carry[19] ,
         \iRF_stage/i_pc_gen/r62/carry[18] ,
         \iRF_stage/i_pc_gen/r62/carry[17] ,
         \iRF_stage/i_pc_gen/r62/carry[16] ,
         \iRF_stage/i_pc_gen/r62/carry[15] ,
         \iRF_stage/i_pc_gen/r62/carry[14] ,
         \iRF_stage/i_pc_gen/r62/carry[13] ,
         \iRF_stage/i_pc_gen/r62/carry[12] ,
         \iRF_stage/i_pc_gen/r62/carry[11] ,
         \iRF_stage/i_pc_gen/r62/carry[10] , \iRF_stage/i_pc_gen/r62/carry[9] ,
         \iRF_stage/i_pc_gen/r62/carry[8] , \iRF_stage/i_pc_gen/r62/carry[7] ,
         \iRF_stage/i_pc_gen/r62/carry[6] , \iRF_stage/i_pc_gen/r62/carry[5] ,
         \iRF_stage/i_pc_gen/r62/carry[4] ,
         \iRF_stage/i_pc_gen/add_70/carry[31] ,
         \iRF_stage/i_pc_gen/add_70/carry[30] ,
         \iRF_stage/i_pc_gen/add_70/carry[29] ,
         \iRF_stage/i_pc_gen/add_70/carry[28] ,
         \iRF_stage/i_pc_gen/add_70/carry[27] ,
         \iRF_stage/i_pc_gen/add_70/carry[26] ,
         \iRF_stage/i_pc_gen/add_70/carry[25] ,
         \iRF_stage/i_pc_gen/add_70/carry[24] ,
         \iRF_stage/i_pc_gen/add_70/carry[23] ,
         \iRF_stage/i_pc_gen/add_70/carry[22] ,
         \iRF_stage/i_pc_gen/add_70/carry[21] ,
         \iRF_stage/i_pc_gen/add_70/carry[20] ,
         \iRF_stage/i_pc_gen/add_70/carry[19] ,
         \iRF_stage/i_pc_gen/add_70/carry[18] ,
         \iRF_stage/i_pc_gen/add_70/carry[17] ,
         \iRF_stage/i_pc_gen/add_70/carry[16] ,
         \iRF_stage/i_pc_gen/add_70/carry[15] ,
         \iRF_stage/i_pc_gen/add_70/carry[14] ,
         \iRF_stage/i_pc_gen/add_70/carry[13] ,
         \iRF_stage/i_pc_gen/add_70/carry[12] ,
         \iRF_stage/i_pc_gen/add_70/carry[11] ,
         \iRF_stage/i_pc_gen/add_70/carry[10] ,
         \iRF_stage/i_pc_gen/add_70/carry[9] ,
         \iRF_stage/i_pc_gen/add_70/carry[8] ,
         \iRF_stage/i_pc_gen/add_70/carry[7] ,
         \iRF_stage/i_pc_gen/add_70/carry[6] ,
         \iRF_stage/i_pc_gen/add_70/carry[5] ,
         \iRF_stage/i_pc_gen/add_70/carry[4] ,
         \iRF_stage/i_pc_gen/add_70/carry[3] ,
         \iRF_stage/i_pc_gen/add_70/carry[2] ,
         \iRF_stage/i_pc_gen/add_70/carry[1] ,
         \iRF_stage/MAIN_FSM/add_58/carry[5] ,
         \iRF_stage/MAIN_FSM/add_58/carry[4] ,
         \iRF_stage/MAIN_FSM/add_58/carry[3] ,
         \iRF_stage/MAIN_FSM/add_58/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n302, n303, n304, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939;
  wire   [31:0] BUS9884;
  wire   [3:0] BUS5985;
  wire   [31:0] BUS22401;
  wire   [31:0] BUS7219;
  wire   [31:0] BUS15471;
  wire   [31:0] BUS27031;
  wire   [4:0] BUS775;
  wire   [4:0] BUS748;
  wire   [31:0] BUS24839;
  wire   [4:0] BUS756;
  wire   [31:0] BUS7160;
  wire   [4:0] BUS18211;
  wire   [31:0] BUS7231;
  wire   [31:0] BUS7101;
  wire   [31:0] BUS7117;
  wire   [31:0] BUS422;
  wire   [31:0] BUS7772;
  wire   [4:0] BUS1724;
  wire   [4:0] BUS1726;
  assign \iRF_stage/BUS3236[4]  = ins_i[20];
  assign \iRF_stage/BUS3236[3]  = ins_i[19];
  assign \iRF_stage/BUS3236[2]  = ins_i[18];
  assign \iRF_stage/BUS3236[1]  = ins_i[17];
  assign \iRF_stage/BUS3236[0]  = ins_i[16];
  assign \iRF_stage/BUS3237[4]  = ins_i[25];
  assign \iRF_stage/BUS3237[3]  = ins_i[24];
  assign \iRF_stage/BUS3237[2]  = ins_i[23];
  assign \iRF_stage/BUS3237[1]  = ins_i[22];
  assign \iRF_stage/BUS3237[0]  = ins_i[21];

  EDFFX4 \iRF_stage/reg_bank/r_rdaddress_b_reg_3_  ( .D(\iRF_stage/BUS3236[3] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N20 ), .QN(n342) );
  EDFFX4 \iRF_stage/reg_bank/r_rdaddress_a_reg_3_  ( .D(\iRF_stage/BUS3237[3] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N15 ), .QN(n337) );
  EDFFTRX1 \iRF_stage/MAIN_FSM/riack_reg  ( .RN(rst), .D(
        \iRF_stage/MAIN_FSM/CurrState[0] ), .E(n1935), .CK(clk), .QN(n304) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_0_  ( .RN(n1933), .D(ins_i[0]), .E(
        n1936), .CK(clk), .QN(n317) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_1_  ( .RN(n1933), .D(ins_i[1]), .E(
        n1936), .CK(clk), .QN(n326) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_2_  ( .RN(n1933), .D(ins_i[2]), .E(
        n1936), .CK(clk), .QN(n327) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_3_  ( .RN(n1933), .D(ins_i[3]), .E(
        n1936), .CK(clk), .QN(n328) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_4_  ( .RN(n1933), .D(ins_i[4]), .E(
        n1936), .CK(clk), .QN(n329) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_5_  ( .RN(n1933), .D(ins_i[5]), .E(
        n1936), .CK(clk), .QN(n330) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_6_  ( .RN(n1933), .D(ins_i[6]), .E(
        n1936), .CK(clk), .QN(n331) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_7_  ( .RN(n1933), .D(ins_i[7]), .E(
        n1936), .CK(clk), .QN(n332) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_8_  ( .RN(n1933), .D(ins_i[8]), .E(
        n1936), .CK(clk), .QN(n307) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_9_  ( .RN(n1933), .D(ins_i[9]), .E(
        n1936), .CK(clk), .QN(n308) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_10_  ( .RN(n1933), .D(ins_i[10]), .E(
        n1936), .CK(clk), .QN(n309) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_11_  ( .RN(n1933), .D(ins_i[11]), .E(
        n1936), .CK(clk), .QN(n310) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_12_  ( .RN(n1933), .D(ins_i[12]), .E(
        n1936), .CK(clk), .QN(n311) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_13_  ( .RN(n1933), .D(ins_i[13]), .E(
        n1936), .CK(clk), .QN(n312) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_14_  ( .RN(n1933), .D(ins_i[14]), .E(
        n1936), .CK(clk), .QN(n313) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_15_  ( .RN(n1933), .D(ins_i[15]), .E(
        n1936), .CK(clk), .Q(n44), .QN(n314) );
  EDFFTRX1 \decoder_pipe/pipereg/U2/cmp_ctl_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2056[0] ), .E(n1936), .CK(clk), .QN(n293) );
  EDFFTRX1 \decoder_pipe/pipereg/U2/cmp_ctl_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2056[1] ), .E(n1936), .CK(clk), .QN(n294) );
  EDFFTRX1 \decoder_pipe/pipereg/U2/cmp_ctl_o_reg_2_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2056[2] ), .E(n1936), .CK(clk), .QN(n295) );
  EDFFTRX1 \decoder_pipe/pipereg/U4/ext_ctl_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2072[0] ), .E(n1936), .CK(clk), .QN(n296) );
  EDFFTRX1 \decoder_pipe/pipereg/U4/ext_ctl_o_reg_1_  ( .RN(n1933), .D(n1930), 
        .E(n1936), .CK(clk), .QN(n297) );
  EDFFTRX1 \decoder_pipe/pipereg/U4/ext_ctl_o_reg_2_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2072[2] ), .E(n1936), .CK(clk), .Q(n42), .QN(n298) );
  EDFFTRX1 \decoder_pipe/pipereg/U5/rd_sel_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2110[0] ), .E(n1936), .CK(clk), .QN(n299) );
  EDFFTRX1 \decoder_pipe/pipereg/U5/rd_sel_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2110[1] ), .E(n1936), .CK(clk), .QN(n300) );
  EDFFTRX1 \decoder_pipe/pipereg/U8/pc_gen_ctl_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2102[0] ), .E(n1936), .CK(clk), .Q(n38) );
  EDFFTRX1 \decoder_pipe/pipereg/U8/pc_gen_ctl_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2102[1] ), .E(n1936), .CK(clk), .QN(n302) );
  EDFFTRX1 \decoder_pipe/pipereg/U8/pc_gen_ctl_o_reg_2_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2102[2] ), .E(n1936), .CK(clk), .QN(n303) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_0_  ( .D(\iRF_stage/i_pc_gen/N34 ), .E(
        n1932), .CK(clk), .Q(n76) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_1_  ( .D(BUS27031[1]), .E(n1932), .CK(clk), 
        .Q(n75) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_2_  ( .D(BUS27031[2]), .E(n1932), .CK(clk), 
        .Q(n69) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_3_  ( .D(BUS27031[3]), .E(n1932), .CK(clk), 
        .Q(n68) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_4_  ( .D(BUS27031[4]), .E(n1932), .CK(clk), 
        .Q(n70) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_5_  ( .D(BUS27031[5]), .E(n1932), .CK(clk), 
        .Q(n57) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_6_  ( .D(BUS27031[6]), .E(n1932), .CK(clk), 
        .Q(n56) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_7_  ( .D(BUS27031[7]), .E(n1932), .CK(clk), 
        .Q(n55) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_8_  ( .D(BUS27031[8]), .E(n1932), .CK(clk), 
        .Q(n58) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_9_  ( .D(BUS27031[9]), .E(n1932), .CK(clk), 
        .Q(n54) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_10_  ( .D(BUS27031[10]), .E(n1932), .CK(
        clk), .Q(n59) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_11_  ( .D(BUS27031[11]), .E(n1932), .CK(
        clk), .Q(n60) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_12_  ( .D(BUS27031[12]), .E(n1932), .CK(
        clk), .Q(n53) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_13_  ( .D(BUS27031[13]), .E(n1932), .CK(
        clk), .Q(n52) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_14_  ( .D(BUS27031[14]), .E(n1932), .CK(
        clk), .Q(n61) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_15_  ( .D(BUS27031[15]), .E(n1932), .CK(
        clk), .Q(n51) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_16_  ( .D(BUS27031[16]), .E(n1932), .CK(
        clk), .Q(n62) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_17_  ( .D(BUS27031[17]), .E(n1932), .CK(
        clk), .Q(n63) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_18_  ( .D(BUS27031[18]), .E(n1932), .CK(
        clk), .Q(n50) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_19_  ( .D(BUS27031[19]), .E(n1932), .CK(
        clk), .Q(n49) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_20_  ( .D(BUS27031[20]), .E(n1932), .CK(
        clk), .Q(n64) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_21_  ( .D(BUS27031[21]), .E(n1932), .CK(
        clk), .Q(n48) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_22_  ( .D(BUS27031[22]), .E(n1932), .CK(
        clk), .Q(n65) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_23_  ( .D(BUS27031[23]), .E(n1932), .CK(
        clk), .Q(n66) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_24_  ( .D(BUS27031[24]), .E(n1932), .CK(
        clk), .Q(n47) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_25_  ( .D(BUS27031[25]), .E(n1932), .CK(
        clk), .Q(n46) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_26_  ( .D(BUS27031[26]), .E(n1932), .CK(
        clk), .Q(n67) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_27_  ( .D(BUS27031[27]), .E(n1932), .CK(
        clk), .Q(n45) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_28_  ( .D(BUS27031[28]), .E(n1932), .CK(
        clk), .Q(n73) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_29_  ( .D(BUS27031[29]), .E(n1932), .CK(
        clk), .Q(n72) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_30_  ( .D(BUS27031[30]), .E(n1932), .CK(
        clk), .Q(n71) );
  EDFFX1 \iexec_stage/spc/r32_o_reg_31_  ( .D(BUS27031[31]), .E(n1932), .CK(
        clk), .Q(n74) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_0_  ( .D(BUS15471[0]), .CK(clk), .Q(n34) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_1_  ( .D(BUS15471[1]), .CK(clk), .Q(n23) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_2_  ( .D(BUS15471[2]), .CK(clk), .Q(n12) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_3_  ( .D(BUS15471[3]), .CK(clk), .Q(n9)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_4_  ( .D(BUS15471[4]), .CK(clk), .Q(n8)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_5_  ( .D(BUS15471[5]), .CK(clk), .Q(n7)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_6_  ( .D(BUS15471[6]), .CK(clk), .Q(n6)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_7_  ( .D(BUS15471[7]), .CK(clk), .Q(n5)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_8_  ( .D(BUS15471[8]), .CK(clk), .Q(n4)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_9_  ( .D(BUS15471[9]), .CK(clk), .Q(n3)
         );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_10_  ( .D(BUS15471[10]), .CK(clk), .Q(
        n33) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_11_  ( .D(BUS15471[11]), .CK(clk), .Q(
        n32) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_12_  ( .D(BUS15471[12]), .CK(clk), .Q(
        n31) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_13_  ( .D(BUS15471[13]), .CK(clk), .Q(
        n30) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_14_  ( .D(BUS15471[14]), .CK(clk), .Q(
        n29) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_15_  ( .D(BUS15471[15]), .CK(clk), .Q(
        n28) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_16_  ( .D(BUS15471[16]), .CK(clk), .Q(
        n27) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_17_  ( .D(BUS15471[17]), .CK(clk), .Q(
        n26) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_18_  ( .D(BUS15471[18]), .CK(clk), .Q(
        n25) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_19_  ( .D(BUS15471[19]), .CK(clk), .Q(
        n24) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_20_  ( .D(BUS15471[20]), .CK(clk), .Q(
        n22) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_21_  ( .D(BUS15471[21]), .CK(clk), .Q(
        n21) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_22_  ( .D(BUS15471[22]), .CK(clk), .Q(
        n20) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_23_  ( .D(BUS15471[23]), .CK(clk), .Q(
        n19) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_24_  ( .D(BUS15471[24]), .CK(clk), .Q(
        n18) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_25_  ( .D(BUS15471[25]), .CK(clk), .Q(
        n17) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_26_  ( .D(BUS15471[26]), .CK(clk), .Q(
        n16) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_27_  ( .D(BUS15471[27]), .CK(clk), .Q(
        n15) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_28_  ( .D(BUS15471[28]), .CK(clk), .Q(
        n14) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_29_  ( .D(BUS15471[29]), .CK(clk), .Q(
        n13) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_30_  ( .D(BUS15471[30]), .CK(clk), .Q(
        n11) );
  DFFX1 \iRF_stage/reg_bank/r_data_reg_31_  ( .D(BUS15471[31]), .CK(clk), .Q(
        n10) );
  DFFTRX1 \MEM_CTL/dmem_ctl_post/ctl_o_reg_0_  ( .D(BUS5985[0]), .RN(n1878), 
        .CK(clk), .Q(n35), .QN(n276) );
  DFFTRX1 \MEM_CTL/dmem_ctl_post/ctl_o_reg_1_  ( .D(BUS5985[1]), .RN(n1878), 
        .CK(clk), .QN(n277) );
  DFFTRX1 \MEM_CTL/dmem_ctl_post/ctl_o_reg_2_  ( .D(BUS5985[2]), .RN(n1878), 
        .CK(clk), .Q(n2), .QN(n278) );
  DFFTRX1 \MEM_CTL/dmem_ctl_post/ctl_o_reg_3_  ( .D(BUS5985[3]), .RN(n1878), 
        .CK(clk), .Q(n43), .QN(n279) );
  DFFTRX1 \iRF_stage/MAIN_FSM/CurrState_reg_3_  ( .D(n1929), .RN(rst), .CK(clk), .Q(n37), .QN(\iRF_stage/MAIN_FSM/n17 ) );
  DFFTRX1 \iRF_stage/MAIN_FSM/delay_counter_reg_5_  ( .D(
        \iRF_stage/MAIN_FSM/N37 ), .RN(\iRF_stage/MAIN_FSM/n57 ), .CK(clk), 
        .Q(n41) );
  DFFTRX1 \decoder_pipe/pipereg/U14/muxb_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5483[0] ), .RN(n1934), .CK(clk), .QN(n280) );
  DFFTRX1 \decoder_pipe/pipereg/U14/muxb_ctl_o_reg_1_  ( .D(
        \decoder_pipe/pipereg/BUS5483[1] ), .RN(n1934), .CK(clk), .QN(n281) );
  DFFTRX1 \decoder_pipe/pipereg/U16/alu_func_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5674[0] ), .RN(n1934), .CK(clk), .Q(n40), 
        .QN(n286) );
  DFFTRX1 \decoder_pipe/pipereg/U16/alu_func_o_reg_1_  ( .D(
        \decoder_pipe/pipereg/BUS5674[1] ), .RN(n1934), .CK(clk), .Q(n39), 
        .QN(n287) );
  DFFTRX1 \decoder_pipe/pipereg/U16/alu_func_o_reg_2_  ( .D(
        \decoder_pipe/pipereg/BUS5674[2] ), .RN(n1934), .CK(clk), .QN(n288) );
  DFFTRX1 \decoder_pipe/pipereg/U16/alu_func_o_reg_3_  ( .D(
        \decoder_pipe/pipereg/BUS5674[3] ), .RN(n1934), .CK(clk), .QN(n289) );
  DFFTRX1 \decoder_pipe/pipereg/U16/alu_func_o_reg_4_  ( .D(
        \decoder_pipe/pipereg/BUS5674[4] ), .RN(n1934), .CK(clk), .Q(n36), 
        .QN(n290) );
  DFFTRX1 \decoder_pipe/pipereg/U17/muxa_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5008[0] ), .RN(n1934), .CK(clk), .QN(n291) );
  DFFTRX1 \decoder_pipe/pipereg/U17/muxa_ctl_o_reg_1_  ( .D(
        \decoder_pipe/pipereg/BUS5008[1] ), .RN(n1934), .CK(clk), .Q(n77), 
        .QN(n292) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_0_  ( .D(BUS22401[0]), .CK(clk), .Q(
        BUS7772[0]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_1_  ( .D(BUS22401[1]), .CK(clk), .Q(
        BUS7772[1]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_2_  ( .D(BUS22401[2]), .CK(clk), .Q(
        BUS7772[2]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_3_  ( .D(BUS22401[3]), .CK(clk), .Q(
        BUS7772[3]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_4_  ( .D(BUS22401[4]), .CK(clk), .Q(
        BUS7772[4]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_5_  ( .D(BUS22401[5]), .CK(clk), .Q(
        BUS7772[5]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_6_  ( .D(BUS22401[6]), .CK(clk), .Q(
        BUS7772[6]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_7_  ( .D(BUS22401[7]), .CK(clk), .Q(
        BUS7772[7]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_8_  ( .D(BUS22401[8]), .CK(clk), .Q(
        BUS7772[8]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_9_  ( .D(BUS22401[9]), .CK(clk), .Q(
        BUS7772[9]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_10_  ( .D(BUS22401[10]), .CK(clk), .Q(
        BUS7772[10]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_11_  ( .D(BUS22401[11]), .CK(clk), .Q(
        BUS7772[11]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_12_  ( .D(BUS22401[12]), .CK(clk), .Q(
        BUS7772[12]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_13_  ( .D(BUS22401[13]), .CK(clk), .Q(
        BUS7772[13]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_14_  ( .D(BUS22401[14]), .CK(clk), .Q(
        BUS7772[14]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_15_  ( .D(BUS22401[15]), .CK(clk), .Q(
        BUS7772[15]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_16_  ( .D(BUS22401[16]), .CK(clk), .Q(
        BUS7772[16]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_17_  ( .D(BUS22401[17]), .CK(clk), .Q(
        BUS7772[17]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_18_  ( .D(BUS22401[18]), .CK(clk), .Q(
        BUS7772[18]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_19_  ( .D(BUS22401[19]), .CK(clk), .Q(
        BUS7772[19]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_20_  ( .D(BUS22401[20]), .CK(clk), .Q(
        BUS7772[20]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_21_  ( .D(BUS22401[21]), .CK(clk), .Q(
        BUS7772[21]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_22_  ( .D(BUS22401[22]), .CK(clk), .Q(
        BUS7772[22]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_23_  ( .D(BUS22401[23]), .CK(clk), .Q(
        BUS7772[23]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_24_  ( .D(BUS22401[24]), .CK(clk), .Q(
        BUS7772[24]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_25_  ( .D(BUS22401[25]), .CK(clk), .Q(
        BUS7772[25]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_26_  ( .D(BUS22401[26]), .CK(clk), .Q(
        BUS7772[26]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_27_  ( .D(BUS22401[27]), .CK(clk), .Q(
        BUS7772[27]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_28_  ( .D(BUS22401[28]), .CK(clk), .Q(
        BUS7772[28]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_29_  ( .D(BUS22401[29]), .CK(clk), .Q(
        BUS7772[29]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_30_  ( .D(BUS22401[30]), .CK(clk), .Q(
        BUS7772[30]) );
  DFFHQX1 \cop_dout_reg/r32_o_reg_31_  ( .D(BUS22401[31]), .CK(clk), .Q(
        BUS7772[31]) );
  DFFHQX1 \decoder_pipe/pipereg/U20/wb_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5682[0] ), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS7822[0] ) );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_16_  ( .RN(n1933), .D(
        \iRF_stage/BUS3236[0] ), .E(n1936), .CK(clk), .Q(BUS756[0]), .QN(n315)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_17_  ( .RN(n1933), .D(
        \iRF_stage/BUS3236[1] ), .E(n1936), .CK(clk), .Q(BUS756[1]), .QN(n316)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_18_  ( .RN(n1933), .D(
        \iRF_stage/BUS3236[2] ), .E(n1936), .CK(clk), .Q(BUS756[2]), .QN(n318)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_19_  ( .RN(n1933), .D(
        \iRF_stage/BUS3236[3] ), .E(n1936), .CK(clk), .Q(BUS756[3]), .QN(n319)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_20_  ( .RN(n1933), .D(
        \iRF_stage/BUS3236[4] ), .E(n1936), .CK(clk), .Q(BUS756[4]), .QN(n320)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_21_  ( .RN(n1933), .D(
        \iRF_stage/BUS3237[0] ), .E(n1936), .CK(clk), .Q(BUS748[0]), .QN(n321)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_22_  ( .RN(n1933), .D(
        \iRF_stage/BUS3237[1] ), .E(n1936), .CK(clk), .Q(BUS748[1]), .QN(n322)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_23_  ( .RN(n1933), .D(
        \iRF_stage/BUS3237[2] ), .E(n1936), .CK(clk), .Q(BUS748[2]), .QN(n323)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_24_  ( .RN(n1933), .D(
        \iRF_stage/BUS3237[3] ), .E(n1936), .CK(clk), .Q(BUS748[3]), .QN(n324)
         );
  EDFFTRX1 \iRF_stage/ins_reg/r32_o_reg_25_  ( .RN(n1933), .D(
        \iRF_stage/BUS3237[4] ), .E(n1936), .CK(clk), .Q(BUS748[4]), .QN(n325)
         );
  DFFHQX1 \rt_reg/r32_o_reg_0_  ( .D(BUS7160[0]), .CK(clk), .Q(BUS7117[0]) );
  DFFHQX1 \rt_reg/r32_o_reg_1_  ( .D(BUS7160[1]), .CK(clk), .Q(BUS7117[1]) );
  DFFHQX1 \rt_reg/r32_o_reg_2_  ( .D(BUS7160[2]), .CK(clk), .Q(BUS7117[2]) );
  DFFHQX1 \rt_reg/r32_o_reg_3_  ( .D(BUS7160[3]), .CK(clk), .Q(BUS7117[3]) );
  DFFHQX1 \rt_reg/r32_o_reg_4_  ( .D(BUS7160[4]), .CK(clk), .Q(BUS7117[4]) );
  DFFHQX1 \rt_reg/r32_o_reg_5_  ( .D(BUS7160[5]), .CK(clk), .Q(BUS7117[5]) );
  DFFHQX1 \rt_reg/r32_o_reg_6_  ( .D(BUS7160[6]), .CK(clk), .Q(BUS7117[6]) );
  DFFHQX1 \rt_reg/r32_o_reg_7_  ( .D(BUS7160[7]), .CK(clk), .Q(BUS7117[7]) );
  DFFHQX1 \rt_reg/r32_o_reg_8_  ( .D(BUS7160[8]), .CK(clk), .Q(BUS7117[8]) );
  DFFHQX1 \rt_reg/r32_o_reg_9_  ( .D(BUS7160[9]), .CK(clk), .Q(BUS7117[9]) );
  DFFHQX1 \rt_reg/r32_o_reg_10_  ( .D(BUS7160[10]), .CK(clk), .Q(BUS7117[10])
         );
  DFFHQX1 \rt_reg/r32_o_reg_11_  ( .D(BUS7160[11]), .CK(clk), .Q(BUS7117[11])
         );
  DFFHQX1 \rt_reg/r32_o_reg_12_  ( .D(BUS7160[12]), .CK(clk), .Q(BUS7117[12])
         );
  DFFHQX1 \rt_reg/r32_o_reg_13_  ( .D(BUS7160[13]), .CK(clk), .Q(BUS7117[13])
         );
  DFFHQX1 \rt_reg/r32_o_reg_14_  ( .D(BUS7160[14]), .CK(clk), .Q(BUS7117[14])
         );
  DFFHQX1 \rt_reg/r32_o_reg_15_  ( .D(BUS7160[15]), .CK(clk), .Q(BUS7117[15])
         );
  DFFHQX1 \rt_reg/r32_o_reg_16_  ( .D(BUS7160[16]), .CK(clk), .Q(BUS7117[16])
         );
  DFFHQX1 \rt_reg/r32_o_reg_17_  ( .D(BUS7160[17]), .CK(clk), .Q(BUS7117[17])
         );
  DFFHQX1 \rt_reg/r32_o_reg_18_  ( .D(BUS7160[18]), .CK(clk), .Q(BUS7117[18])
         );
  DFFHQX1 \rt_reg/r32_o_reg_19_  ( .D(BUS7160[19]), .CK(clk), .Q(BUS7117[19])
         );
  DFFHQX1 \rt_reg/r32_o_reg_20_  ( .D(BUS7160[20]), .CK(clk), .Q(BUS7117[20])
         );
  DFFHQX1 \rt_reg/r32_o_reg_21_  ( .D(BUS7160[21]), .CK(clk), .Q(BUS7117[21])
         );
  DFFHQX1 \rt_reg/r32_o_reg_22_  ( .D(BUS7160[22]), .CK(clk), .Q(BUS7117[22])
         );
  DFFHQX1 \rt_reg/r32_o_reg_23_  ( .D(BUS7160[23]), .CK(clk), .Q(BUS7117[23])
         );
  DFFHQX1 \rt_reg/r32_o_reg_24_  ( .D(BUS7160[24]), .CK(clk), .Q(BUS7117[24])
         );
  DFFHQX1 \rt_reg/r32_o_reg_25_  ( .D(BUS7160[25]), .CK(clk), .Q(BUS7117[25])
         );
  DFFHQX1 \rt_reg/r32_o_reg_26_  ( .D(BUS7160[26]), .CK(clk), .Q(BUS7117[26])
         );
  DFFHQX1 \rt_reg/r32_o_reg_27_  ( .D(BUS7160[27]), .CK(clk), .Q(BUS7117[27])
         );
  DFFHQX1 \rt_reg/r32_o_reg_28_  ( .D(BUS7160[28]), .CK(clk), .Q(BUS7117[28])
         );
  DFFHQX1 \rt_reg/r32_o_reg_29_  ( .D(BUS7160[29]), .CK(clk), .Q(BUS7117[29])
         );
  DFFHQX1 \rt_reg/r32_o_reg_30_  ( .D(BUS7160[30]), .CK(clk), .Q(BUS7117[30])
         );
  DFFHQX1 \rt_reg/r32_o_reg_31_  ( .D(BUS7160[31]), .CK(clk), .Q(BUS7117[31])
         );
  DFFHQX1 \rs_reg/r32_o_reg_0_  ( .D(BUS24839[0]), .CK(clk), .Q(BUS7101[0]) );
  DFFHQX1 \rs_reg/r32_o_reg_1_  ( .D(BUS24839[1]), .CK(clk), .Q(BUS7101[1]) );
  DFFHQX1 \rs_reg/r32_o_reg_2_  ( .D(BUS24839[2]), .CK(clk), .Q(BUS7101[2]) );
  DFFHQX1 \rs_reg/r32_o_reg_3_  ( .D(BUS24839[3]), .CK(clk), .Q(BUS7101[3]) );
  DFFHQX1 \rs_reg/r32_o_reg_4_  ( .D(BUS24839[4]), .CK(clk), .Q(BUS7101[4]) );
  DFFHQX1 \rs_reg/r32_o_reg_5_  ( .D(BUS24839[5]), .CK(clk), .Q(BUS7101[5]) );
  DFFHQX1 \rs_reg/r32_o_reg_6_  ( .D(BUS24839[6]), .CK(clk), .Q(BUS7101[6]) );
  DFFHQX1 \rs_reg/r32_o_reg_7_  ( .D(BUS24839[7]), .CK(clk), .Q(BUS7101[7]) );
  DFFHQX1 \rs_reg/r32_o_reg_8_  ( .D(BUS24839[8]), .CK(clk), .Q(BUS7101[8]) );
  DFFHQX1 \rs_reg/r32_o_reg_9_  ( .D(BUS24839[9]), .CK(clk), .Q(BUS7101[9]) );
  DFFHQX1 \rs_reg/r32_o_reg_10_  ( .D(BUS24839[10]), .CK(clk), .Q(BUS7101[10])
         );
  DFFHQX1 \rs_reg/r32_o_reg_11_  ( .D(BUS24839[11]), .CK(clk), .Q(BUS7101[11])
         );
  DFFHQX1 \rs_reg/r32_o_reg_12_  ( .D(BUS24839[12]), .CK(clk), .Q(BUS7101[12])
         );
  DFFHQX1 \rs_reg/r32_o_reg_13_  ( .D(BUS24839[13]), .CK(clk), .Q(BUS7101[13])
         );
  DFFHQX1 \rs_reg/r32_o_reg_14_  ( .D(BUS24839[14]), .CK(clk), .Q(BUS7101[14])
         );
  DFFHQX1 \rs_reg/r32_o_reg_15_  ( .D(BUS24839[15]), .CK(clk), .Q(BUS7101[15])
         );
  DFFHQX1 \rs_reg/r32_o_reg_16_  ( .D(BUS24839[16]), .CK(clk), .Q(BUS7101[16])
         );
  DFFHQX1 \rs_reg/r32_o_reg_17_  ( .D(BUS24839[17]), .CK(clk), .Q(BUS7101[17])
         );
  DFFHQX1 \rs_reg/r32_o_reg_18_  ( .D(BUS24839[18]), .CK(clk), .Q(BUS7101[18])
         );
  DFFHQX1 \rs_reg/r32_o_reg_19_  ( .D(BUS24839[19]), .CK(clk), .Q(BUS7101[19])
         );
  DFFHQX1 \rs_reg/r32_o_reg_20_  ( .D(BUS24839[20]), .CK(clk), .Q(BUS7101[20])
         );
  DFFHQX1 \rs_reg/r32_o_reg_21_  ( .D(BUS24839[21]), .CK(clk), .Q(BUS7101[21])
         );
  DFFHQX1 \rs_reg/r32_o_reg_22_  ( .D(BUS24839[22]), .CK(clk), .Q(BUS7101[22])
         );
  DFFHQX1 \rs_reg/r32_o_reg_23_  ( .D(BUS24839[23]), .CK(clk), .Q(BUS7101[23])
         );
  DFFHQX1 \rs_reg/r32_o_reg_24_  ( .D(BUS24839[24]), .CK(clk), .Q(BUS7101[24])
         );
  DFFHQX1 \rs_reg/r32_o_reg_25_  ( .D(BUS24839[25]), .CK(clk), .Q(BUS7101[25])
         );
  DFFHQX1 \rs_reg/r32_o_reg_26_  ( .D(BUS24839[26]), .CK(clk), .Q(BUS7101[26])
         );
  DFFHQX1 \rs_reg/r32_o_reg_27_  ( .D(BUS24839[27]), .CK(clk), .Q(BUS7101[27])
         );
  DFFHQX1 \rs_reg/r32_o_reg_28_  ( .D(BUS24839[28]), .CK(clk), .Q(BUS7101[28])
         );
  DFFHQX1 \rs_reg/r32_o_reg_29_  ( .D(BUS24839[29]), .CK(clk), .Q(BUS7101[29])
         );
  DFFHQX1 \rs_reg/r32_o_reg_30_  ( .D(BUS24839[30]), .CK(clk), .Q(BUS7101[30])
         );
  DFFHQX1 \rs_reg/r32_o_reg_31_  ( .D(BUS24839[31]), .CK(clk), .Q(BUS7101[31])
         );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_0_  ( .D(\iRF_stage/i_pc_gen/N34 ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[0] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_1_  ( .D(BUS27031[1]), .CK(clk), .Q(
        \iexec_stage/BUS2332[1] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_2_  ( .D(n1939), .CK(clk), .Q(
        \iexec_stage/BUS2332[2] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_3_  ( .D(\iexec_stage/BUS2446[3] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[3] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_4_  ( .D(\iexec_stage/BUS2446[4] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[4] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_5_  ( .D(\iexec_stage/BUS2446[5] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[5] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_6_  ( .D(\iexec_stage/BUS2446[6] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[6] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_7_  ( .D(\iexec_stage/BUS2446[7] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[7] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_8_  ( .D(\iexec_stage/BUS2446[8] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[8] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_9_  ( .D(\iexec_stage/BUS2446[9] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[9] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_10_  ( .D(\iexec_stage/BUS2446[10] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[10] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_11_  ( .D(\iexec_stage/BUS2446[11] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[11] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_12_  ( .D(\iexec_stage/BUS2446[12] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[12] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_13_  ( .D(\iexec_stage/BUS2446[13] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[13] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_14_  ( .D(\iexec_stage/BUS2446[14] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[14] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_15_  ( .D(\iexec_stage/BUS2446[15] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[15] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_16_  ( .D(\iexec_stage/BUS2446[16] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[16] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_17_  ( .D(\iexec_stage/BUS2446[17] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[17] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_18_  ( .D(\iexec_stage/BUS2446[18] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[18] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_19_  ( .D(\iexec_stage/BUS2446[19] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[19] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_20_  ( .D(\iexec_stage/BUS2446[20] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[20] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_21_  ( .D(\iexec_stage/BUS2446[21] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[21] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_22_  ( .D(\iexec_stage/BUS2446[22] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[22] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_23_  ( .D(\iexec_stage/BUS2446[23] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[23] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_24_  ( .D(\iexec_stage/BUS2446[24] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[24] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_25_  ( .D(\iexec_stage/BUS2446[25] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[25] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_26_  ( .D(\iexec_stage/BUS2446[26] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[26] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_27_  ( .D(\iexec_stage/BUS2446[27] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[27] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_28_  ( .D(\iexec_stage/BUS2446[28] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[28] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_29_  ( .D(\iexec_stage/BUS2446[29] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[29] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_30_  ( .D(\iexec_stage/BUS2446[30] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[30] ) );
  DFFHQX1 \iexec_stage/pc_nxt/r32_o_reg_31_  ( .D(\iexec_stage/BUS2446[31] ), 
        .CK(clk), .Q(\iexec_stage/BUS2332[31] ) );
  DFFHQX1 \alu_pass1/r32_o_reg_0_  ( .D(cop_addr_o[0]), .CK(clk), .Q(BUS422[0]) );
  DFFHQX1 \alu_pass1/r32_o_reg_1_  ( .D(cop_addr_o[1]), .CK(clk), .Q(BUS422[1]) );
  DFFHQX1 \alu_pass1/r32_o_reg_2_  ( .D(cop_addr_o[2]), .CK(clk), .Q(BUS422[2]) );
  DFFHQX1 \alu_pass1/r32_o_reg_3_  ( .D(cop_addr_o[3]), .CK(clk), .Q(BUS422[3]) );
  DFFHQX1 \alu_pass1/r32_o_reg_4_  ( .D(cop_addr_o[4]), .CK(clk), .Q(BUS422[4]) );
  DFFHQX1 \alu_pass1/r32_o_reg_5_  ( .D(cop_addr_o[5]), .CK(clk), .Q(BUS422[5]) );
  DFFHQX1 \alu_pass1/r32_o_reg_6_  ( .D(cop_addr_o[6]), .CK(clk), .Q(BUS422[6]) );
  DFFHQX1 \alu_pass1/r32_o_reg_7_  ( .D(cop_addr_o[7]), .CK(clk), .Q(BUS422[7]) );
  DFFHQX1 \alu_pass1/r32_o_reg_8_  ( .D(cop_addr_o[8]), .CK(clk), .Q(BUS422[8]) );
  DFFHQX1 \alu_pass1/r32_o_reg_9_  ( .D(cop_addr_o[9]), .CK(clk), .Q(BUS422[9]) );
  DFFHQX1 \alu_pass1/r32_o_reg_10_  ( .D(cop_addr_o[10]), .CK(clk), .Q(
        BUS422[10]) );
  DFFHQX1 \alu_pass1/r32_o_reg_11_  ( .D(cop_addr_o[11]), .CK(clk), .Q(
        BUS422[11]) );
  DFFHQX1 \alu_pass1/r32_o_reg_12_  ( .D(cop_addr_o[12]), .CK(clk), .Q(
        BUS422[12]) );
  DFFHQX1 \alu_pass1/r32_o_reg_13_  ( .D(cop_addr_o[13]), .CK(clk), .Q(
        BUS422[13]) );
  DFFHQX1 \alu_pass1/r32_o_reg_14_  ( .D(cop_addr_o[14]), .CK(clk), .Q(
        BUS422[14]) );
  DFFHQX1 \alu_pass1/r32_o_reg_15_  ( .D(cop_addr_o[15]), .CK(clk), .Q(
        BUS422[15]) );
  DFFHQX1 \alu_pass1/r32_o_reg_16_  ( .D(cop_addr_o[16]), .CK(clk), .Q(
        BUS422[16]) );
  DFFHQX1 \alu_pass1/r32_o_reg_17_  ( .D(cop_addr_o[17]), .CK(clk), .Q(
        BUS422[17]) );
  DFFHQX1 \alu_pass1/r32_o_reg_18_  ( .D(cop_addr_o[18]), .CK(clk), .Q(
        BUS422[18]) );
  DFFHQX1 \alu_pass1/r32_o_reg_19_  ( .D(cop_addr_o[19]), .CK(clk), .Q(
        BUS422[19]) );
  DFFHQX1 \alu_pass1/r32_o_reg_20_  ( .D(cop_addr_o[20]), .CK(clk), .Q(
        BUS422[20]) );
  DFFHQX1 \alu_pass1/r32_o_reg_21_  ( .D(cop_addr_o[21]), .CK(clk), .Q(
        BUS422[21]) );
  DFFHQX1 \alu_pass1/r32_o_reg_22_  ( .D(cop_addr_o[22]), .CK(clk), .Q(
        BUS422[22]) );
  DFFHQX1 \alu_pass1/r32_o_reg_23_  ( .D(cop_addr_o[23]), .CK(clk), .Q(
        BUS422[23]) );
  DFFHQX1 \alu_pass1/r32_o_reg_24_  ( .D(cop_addr_o[24]), .CK(clk), .Q(
        BUS422[24]) );
  DFFHQX1 \alu_pass1/r32_o_reg_25_  ( .D(cop_addr_o[25]), .CK(clk), .Q(
        BUS422[25]) );
  DFFHQX1 \alu_pass1/r32_o_reg_26_  ( .D(cop_addr_o[26]), .CK(clk), .Q(
        BUS422[26]) );
  DFFHQX1 \alu_pass1/r32_o_reg_27_  ( .D(cop_addr_o[27]), .CK(clk), .Q(
        BUS422[27]) );
  DFFHQX1 \alu_pass1/r32_o_reg_28_  ( .D(cop_addr_o[28]), .CK(clk), .Q(
        BUS422[28]) );
  DFFHQX1 \alu_pass1/r32_o_reg_29_  ( .D(cop_addr_o[29]), .CK(clk), .Q(
        BUS422[29]) );
  DFFHQX1 \alu_pass1/r32_o_reg_30_  ( .D(cop_addr_o[30]), .CK(clk), .Q(
        BUS422[30]) );
  DFFHQX1 \alu_pass1/r32_o_reg_31_  ( .D(cop_addr_o[31]), .CK(clk), .Q(
        BUS422[31]) );
  DFFHQX1 \decoder_pipe/pipereg/U10/wb_mux_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/U10/n4 ), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5651[0] ) );
  DFFHQX1 \decoder_pipe/pipereg/U11/wb_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/U11/n4 ), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5639[0] ) );
  DFFHQX1 \decoder_pipe/pipereg/U6/alu_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/U6/n4 ), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS4987[0] ) );
  DFFTRX1 \decoder_pipe/pipereg/U15/dmem_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5666[0] ), .RN(n1934), .CK(clk), .Q(
        BUS5985[0]), .QN(n282) );
  DFFTRX1 \decoder_pipe/pipereg/U15/dmem_ctl_o_reg_1_  ( .D(
        \decoder_pipe/pipereg/BUS5666[1] ), .RN(n1934), .CK(clk), .Q(
        BUS5985[1]), .QN(n283) );
  DFFTRX1 \decoder_pipe/pipereg/U15/dmem_ctl_o_reg_2_  ( .D(
        \decoder_pipe/pipereg/BUS5666[2] ), .RN(n1934), .CK(clk), .Q(
        BUS5985[2]), .QN(n284) );
  DFFTRX1 \decoder_pipe/pipereg/U15/dmem_ctl_o_reg_3_  ( .D(
        \decoder_pipe/pipereg/BUS5666[3] ), .RN(n1934), .CK(clk), .Q(
        BUS5985[3]), .QN(n285) );
  DFFHQX1 \decoder_pipe/pipereg/U22/wb_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS7299[0] ), .CK(clk), .Q(NET767) );
  DFFHQX1 \ext_reg/r32_o_reg_1_  ( .D(BUS7219[1]), .CK(clk), .Q(BUS7231[1]) );
  DFFHQX1 \ext_reg/r32_o_reg_2_  ( .D(BUS7219[2]), .CK(clk), .Q(BUS7231[2]) );
  DFFHQX1 \ext_reg/r32_o_reg_3_  ( .D(BUS7219[3]), .CK(clk), .Q(BUS7231[3]) );
  DFFHQX1 \ext_reg/r32_o_reg_4_  ( .D(BUS7219[4]), .CK(clk), .Q(BUS7231[4]) );
  DFFHQX1 \ext_reg/r32_o_reg_5_  ( .D(BUS7219[5]), .CK(clk), .Q(BUS7231[5]) );
  DFFHQX1 \ext_reg/r32_o_reg_6_  ( .D(BUS7219[6]), .CK(clk), .Q(BUS7231[6]) );
  DFFHQX1 \ext_reg/r32_o_reg_7_  ( .D(BUS7219[7]), .CK(clk), .Q(BUS7231[7]) );
  DFFHQX1 \ext_reg/r32_o_reg_8_  ( .D(BUS7219[8]), .CK(clk), .Q(BUS7231[8]) );
  DFFHQX1 \ext_reg/r32_o_reg_9_  ( .D(BUS7219[9]), .CK(clk), .Q(BUS7231[9]) );
  DFFHQX1 \ext_reg/r32_o_reg_10_  ( .D(BUS7219[10]), .CK(clk), .Q(BUS7231[10])
         );
  DFFHQX1 \ext_reg/r32_o_reg_11_  ( .D(BUS7219[11]), .CK(clk), .Q(BUS7231[11])
         );
  DFFHQX1 \ext_reg/r32_o_reg_12_  ( .D(BUS7219[12]), .CK(clk), .Q(BUS7231[12])
         );
  DFFHQX1 \ext_reg/r32_o_reg_13_  ( .D(BUS7219[13]), .CK(clk), .Q(BUS7231[13])
         );
  DFFHQX1 \ext_reg/r32_o_reg_14_  ( .D(BUS7219[14]), .CK(clk), .Q(BUS7231[14])
         );
  DFFHQX1 \ext_reg/r32_o_reg_15_  ( .D(BUS7219[15]), .CK(clk), .Q(BUS7231[15])
         );
  DFFHQX1 \ext_reg/r32_o_reg_16_  ( .D(BUS7219[16]), .CK(clk), .Q(BUS7231[16])
         );
  DFFHQX1 \ext_reg/r32_o_reg_17_  ( .D(BUS7219[17]), .CK(clk), .Q(BUS7231[17])
         );
  DFFHQX1 \ext_reg/r32_o_reg_18_  ( .D(BUS7219[18]), .CK(clk), .Q(BUS7231[18])
         );
  DFFHQX1 \ext_reg/r32_o_reg_19_  ( .D(BUS7219[19]), .CK(clk), .Q(BUS7231[19])
         );
  DFFHQX1 \ext_reg/r32_o_reg_20_  ( .D(BUS7219[20]), .CK(clk), .Q(BUS7231[20])
         );
  DFFHQX1 \ext_reg/r32_o_reg_21_  ( .D(BUS7219[21]), .CK(clk), .Q(BUS7231[21])
         );
  DFFHQX1 \ext_reg/r32_o_reg_22_  ( .D(BUS7219[22]), .CK(clk), .Q(BUS7231[22])
         );
  DFFHQX1 \ext_reg/r32_o_reg_23_  ( .D(BUS7219[23]), .CK(clk), .Q(BUS7231[23])
         );
  DFFHQX1 \ext_reg/r32_o_reg_24_  ( .D(BUS7219[24]), .CK(clk), .Q(BUS7231[24])
         );
  DFFHQX1 \ext_reg/r32_o_reg_25_  ( .D(BUS7219[25]), .CK(clk), .Q(BUS7231[25])
         );
  DFFHQX1 \ext_reg/r32_o_reg_26_  ( .D(BUS7219[26]), .CK(clk), .Q(BUS7231[26])
         );
  DFFHQX1 \ext_reg/r32_o_reg_27_  ( .D(BUS7219[27]), .CK(clk), .Q(BUS7231[27])
         );
  DFFHQX1 \ext_reg/r32_o_reg_28_  ( .D(BUS7219[28]), .CK(clk), .Q(BUS7231[28])
         );
  DFFHQX1 \ext_reg/r32_o_reg_29_  ( .D(BUS7219[29]), .CK(clk), .Q(BUS7231[29])
         );
  DFFHQX1 \ext_reg/r32_o_reg_30_  ( .D(BUS7219[30]), .CK(clk), .Q(BUS7231[30])
         );
  DFFHQX1 \ext_reg/r32_o_reg_31_  ( .D(BUS7219[31]), .CK(clk), .Q(BUS7231[31])
         );
  DFFHQX1 \ext_reg/r32_o_reg_0_  ( .D(BUS7219[0]), .CK(clk), .Q(BUS7231[0]) );
  DFFHQX1 \decoder_pipe/pipereg/U12/wb_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/NET7643 ), .CK(clk), .Q(NET1375) );
  DFFHQX1 \rnd_pass1/r5_o_reg_0_  ( .D(BUS1726[0]), .CK(clk), .Q(BUS1724[0])
         );
  DFFHQX1 \rnd_pass1/r5_o_reg_1_  ( .D(BUS1726[1]), .CK(clk), .Q(BUS1724[1])
         );
  DFFHQX1 \iforward/fw_reg_rns/q_reg_0_  ( .D(BUS748[0]), .CK(clk), .Q(
        \iforward/BUS82[0] ) );
  DFFHQX1 \iforward/fw_reg_rns/q_reg_1_  ( .D(BUS748[1]), .CK(clk), .Q(
        \iforward/BUS82[1] ) );
  DFFHQX1 \iforward/fw_reg_rns/q_reg_2_  ( .D(BUS748[2]), .CK(clk), .Q(
        \iforward/BUS82[2] ) );
  DFFHQX1 \iforward/fw_reg_rns/q_reg_3_  ( .D(BUS748[3]), .CK(clk), .Q(
        \iforward/BUS82[3] ) );
  DFFHQX1 \iforward/fw_reg_rns/q_reg_4_  ( .D(BUS748[4]), .CK(clk), .Q(
        \iforward/BUS82[4] ) );
  DFFHQX1 \iforward/fw_reg_rnt/q_reg_0_  ( .D(BUS756[0]), .CK(clk), .Q(
        \iforward/BUS937[0] ) );
  DFFHQX1 \iforward/fw_reg_rnt/q_reg_1_  ( .D(BUS756[1]), .CK(clk), .Q(
        \iforward/BUS937[1] ) );
  DFFHQX1 \iforward/fw_reg_rnt/q_reg_2_  ( .D(BUS756[2]), .CK(clk), .Q(
        \iforward/BUS937[2] ) );
  DFFHQX1 \iforward/fw_reg_rnt/q_reg_3_  ( .D(BUS756[3]), .CK(clk), .Q(
        \iforward/BUS937[3] ) );
  DFFHQX1 \iforward/fw_reg_rnt/q_reg_4_  ( .D(BUS756[4]), .CK(clk), .Q(
        \iforward/BUS937[4] ) );
  DFFHQX1 \iRF_stage/reg_bank/r_wraddress_reg_4_  ( .D(BUS18211[4]), .CK(clk), 
        .Q(\iRF_stage/reg_bank/r_wraddress[4] ) );
  DFFHQX1 \rnd_pass2/r5_o_reg_4_  ( .D(BUS1724[4]), .CK(clk), .Q(BUS18211[4])
         );
  DFFHQX1 \MEM_CTL/dmem_ctl_post/byte_addr_o_reg_0_  ( .D(addr_o[0]), .CK(clk), 
        .Q(\MEM_CTL/BUS629[0] ) );
  DFFHQX1 \alu_pass0/r32_o_reg_1_  ( .D(addr_o[1]), .CK(clk), .Q(cop_addr_o[1]) );
  DFFHQX1 \alu_pass0/r32_o_reg_2_  ( .D(addr_o[2]), .CK(clk), .Q(cop_addr_o[2]) );
  DFFHQX1 \alu_pass0/r32_o_reg_3_  ( .D(addr_o[3]), .CK(clk), .Q(cop_addr_o[3]) );
  DFFHQX1 \alu_pass0/r32_o_reg_4_  ( .D(addr_o[4]), .CK(clk), .Q(cop_addr_o[4]) );
  DFFHQX1 \alu_pass0/r32_o_reg_5_  ( .D(addr_o[5]), .CK(clk), .Q(cop_addr_o[5]) );
  DFFHQX1 \alu_pass0/r32_o_reg_6_  ( .D(addr_o[6]), .CK(clk), .Q(cop_addr_o[6]) );
  DFFHQX1 \alu_pass0/r32_o_reg_7_  ( .D(addr_o[7]), .CK(clk), .Q(cop_addr_o[7]) );
  DFFHQX1 \alu_pass0/r32_o_reg_8_  ( .D(addr_o[8]), .CK(clk), .Q(cop_addr_o[8]) );
  DFFHQX1 \alu_pass0/r32_o_reg_9_  ( .D(addr_o[9]), .CK(clk), .Q(cop_addr_o[9]) );
  DFFHQX1 \alu_pass0/r32_o_reg_10_  ( .D(addr_o[10]), .CK(clk), .Q(
        cop_addr_o[10]) );
  DFFHQX1 \alu_pass0/r32_o_reg_11_  ( .D(addr_o[11]), .CK(clk), .Q(
        cop_addr_o[11]) );
  DFFHQX1 \alu_pass0/r32_o_reg_12_  ( .D(addr_o[12]), .CK(clk), .Q(
        cop_addr_o[12]) );
  DFFHQX1 \alu_pass0/r32_o_reg_13_  ( .D(addr_o[13]), .CK(clk), .Q(
        cop_addr_o[13]) );
  DFFHQX1 \alu_pass0/r32_o_reg_14_  ( .D(addr_o[14]), .CK(clk), .Q(
        cop_addr_o[14]) );
  DFFHQX1 \alu_pass0/r32_o_reg_15_  ( .D(addr_o[15]), .CK(clk), .Q(
        cop_addr_o[15]) );
  DFFHQX1 \alu_pass0/r32_o_reg_16_  ( .D(addr_o[16]), .CK(clk), .Q(
        cop_addr_o[16]) );
  DFFHQX1 \alu_pass0/r32_o_reg_17_  ( .D(addr_o[17]), .CK(clk), .Q(
        cop_addr_o[17]) );
  DFFHQX1 \alu_pass0/r32_o_reg_18_  ( .D(addr_o[18]), .CK(clk), .Q(
        cop_addr_o[18]) );
  DFFHQX1 \alu_pass0/r32_o_reg_19_  ( .D(addr_o[19]), .CK(clk), .Q(
        cop_addr_o[19]) );
  DFFHQX1 \alu_pass0/r32_o_reg_20_  ( .D(addr_o[20]), .CK(clk), .Q(
        cop_addr_o[20]) );
  DFFHQX1 \alu_pass0/r32_o_reg_21_  ( .D(addr_o[21]), .CK(clk), .Q(
        cop_addr_o[21]) );
  DFFHQX1 \alu_pass0/r32_o_reg_22_  ( .D(addr_o[22]), .CK(clk), .Q(
        cop_addr_o[22]) );
  DFFHQX1 \alu_pass0/r32_o_reg_23_  ( .D(addr_o[23]), .CK(clk), .Q(
        cop_addr_o[23]) );
  DFFHQX1 \alu_pass0/r32_o_reg_24_  ( .D(addr_o[24]), .CK(clk), .Q(
        cop_addr_o[24]) );
  DFFHQX1 \alu_pass0/r32_o_reg_25_  ( .D(addr_o[25]), .CK(clk), .Q(
        cop_addr_o[25]) );
  DFFHQX1 \alu_pass0/r32_o_reg_26_  ( .D(addr_o[26]), .CK(clk), .Q(
        cop_addr_o[26]) );
  DFFHQX1 \alu_pass0/r32_o_reg_27_  ( .D(addr_o[27]), .CK(clk), .Q(
        cop_addr_o[27]) );
  DFFHQX1 \alu_pass0/r32_o_reg_28_  ( .D(addr_o[28]), .CK(clk), .Q(
        cop_addr_o[28]) );
  DFFHQX1 \alu_pass0/r32_o_reg_29_  ( .D(addr_o[29]), .CK(clk), .Q(
        cop_addr_o[29]) );
  DFFHQX1 \alu_pass0/r32_o_reg_30_  ( .D(addr_o[30]), .CK(clk), .Q(
        cop_addr_o[30]) );
  DFFHQX1 \alu_pass0/r32_o_reg_31_  ( .D(addr_o[31]), .CK(clk), .Q(
        cop_addr_o[31]) );
  DFFHQX1 \alu_pass0/r32_o_reg_0_  ( .D(addr_o[0]), .CK(clk), .Q(cop_addr_o[0]) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__0_  ( .D(
        \iRF_stage/reg_bank/n202 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[64] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__1_  ( .D(
        \iRF_stage/reg_bank/n203 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[65] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__2_  ( .D(
        \iRF_stage/reg_bank/n204 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[66] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__3_  ( .D(
        \iRF_stage/reg_bank/n205 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[67] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__4_  ( .D(
        \iRF_stage/reg_bank/n206 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[68] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__5_  ( .D(
        \iRF_stage/reg_bank/n207 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[69] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__6_  ( .D(
        \iRF_stage/reg_bank/n208 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[70] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__7_  ( .D(
        \iRF_stage/reg_bank/n209 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[71] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__8_  ( .D(
        \iRF_stage/reg_bank/n210 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[72] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__9_  ( .D(
        \iRF_stage/reg_bank/n211 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[73] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__10_  ( .D(
        \iRF_stage/reg_bank/n212 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[74] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__11_  ( .D(
        \iRF_stage/reg_bank/n213 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[75] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__12_  ( .D(
        \iRF_stage/reg_bank/n214 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[76] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__13_  ( .D(
        \iRF_stage/reg_bank/n215 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[77] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__14_  ( .D(
        \iRF_stage/reg_bank/n216 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[78] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__15_  ( .D(
        \iRF_stage/reg_bank/n217 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[79] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__16_  ( .D(
        \iRF_stage/reg_bank/n218 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[80] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__17_  ( .D(
        \iRF_stage/reg_bank/n219 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[81] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__18_  ( .D(
        \iRF_stage/reg_bank/n220 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[82] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__19_  ( .D(
        \iRF_stage/reg_bank/n221 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[83] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__20_  ( .D(
        \iRF_stage/reg_bank/n222 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[84] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__21_  ( .D(
        \iRF_stage/reg_bank/n223 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[85] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__22_  ( .D(
        \iRF_stage/reg_bank/n224 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[86] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__23_  ( .D(
        \iRF_stage/reg_bank/n225 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[87] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__24_  ( .D(
        \iRF_stage/reg_bank/n226 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[88] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__25_  ( .D(
        \iRF_stage/reg_bank/n227 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[89] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__26_  ( .D(
        \iRF_stage/reg_bank/n228 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[90] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__27_  ( .D(
        \iRF_stage/reg_bank/n229 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[91] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__28_  ( .D(
        \iRF_stage/reg_bank/n230 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[92] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__29_  ( .D(
        \iRF_stage/reg_bank/n231 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[93] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__30_  ( .D(
        \iRF_stage/reg_bank/n232 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[94] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_29__31_  ( .D(
        \iRF_stage/reg_bank/n233 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[95] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__0_  ( .D(
        \iRF_stage/reg_bank/n330 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[192] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__1_  ( .D(
        \iRF_stage/reg_bank/n331 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[193] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__2_  ( .D(
        \iRF_stage/reg_bank/n332 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[194] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__3_  ( .D(
        \iRF_stage/reg_bank/n333 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[195] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__4_  ( .D(
        \iRF_stage/reg_bank/n334 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[196] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__5_  ( .D(
        \iRF_stage/reg_bank/n335 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[197] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__6_  ( .D(
        \iRF_stage/reg_bank/n336 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[198] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__7_  ( .D(
        \iRF_stage/reg_bank/n337 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[199] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__8_  ( .D(
        \iRF_stage/reg_bank/n338 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[200] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__9_  ( .D(
        \iRF_stage/reg_bank/n339 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[201] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__10_  ( .D(
        \iRF_stage/reg_bank/n340 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[202] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__11_  ( .D(
        \iRF_stage/reg_bank/n341 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[203] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__12_  ( .D(
        \iRF_stage/reg_bank/n342 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[204] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__13_  ( .D(
        \iRF_stage/reg_bank/n343 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[205] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__14_  ( .D(
        \iRF_stage/reg_bank/n344 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[206] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__15_  ( .D(
        \iRF_stage/reg_bank/n345 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[207] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__16_  ( .D(
        \iRF_stage/reg_bank/n346 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[208] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__17_  ( .D(
        \iRF_stage/reg_bank/n347 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[209] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__18_  ( .D(
        \iRF_stage/reg_bank/n348 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[210] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__19_  ( .D(
        \iRF_stage/reg_bank/n349 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[211] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__20_  ( .D(
        \iRF_stage/reg_bank/n350 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[212] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__21_  ( .D(
        \iRF_stage/reg_bank/n351 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[213] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__22_  ( .D(
        \iRF_stage/reg_bank/n352 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[214] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__23_  ( .D(
        \iRF_stage/reg_bank/n353 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[215] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__24_  ( .D(
        \iRF_stage/reg_bank/n354 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[216] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__25_  ( .D(
        \iRF_stage/reg_bank/n355 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[217] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__26_  ( .D(
        \iRF_stage/reg_bank/n356 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[218] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__27_  ( .D(
        \iRF_stage/reg_bank/n357 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[219] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__28_  ( .D(
        \iRF_stage/reg_bank/n358 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[220] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__29_  ( .D(
        \iRF_stage/reg_bank/n359 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[221] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__30_  ( .D(
        \iRF_stage/reg_bank/n360 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[222] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_25__31_  ( .D(
        \iRF_stage/reg_bank/n361 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[223] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__0_  ( .D(
        \iRF_stage/reg_bank/n458 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[320] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__1_  ( .D(
        \iRF_stage/reg_bank/n459 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[321] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__2_  ( .D(
        \iRF_stage/reg_bank/n460 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[322] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__3_  ( .D(
        \iRF_stage/reg_bank/n461 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[323] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__4_  ( .D(
        \iRF_stage/reg_bank/n462 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[324] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__5_  ( .D(
        \iRF_stage/reg_bank/n463 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[325] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__6_  ( .D(
        \iRF_stage/reg_bank/n464 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[326] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__7_  ( .D(
        \iRF_stage/reg_bank/n465 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[327] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__8_  ( .D(
        \iRF_stage/reg_bank/n466 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[328] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__9_  ( .D(
        \iRF_stage/reg_bank/n467 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[329] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__10_  ( .D(
        \iRF_stage/reg_bank/n468 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[330] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__11_  ( .D(
        \iRF_stage/reg_bank/n469 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[331] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__12_  ( .D(
        \iRF_stage/reg_bank/n470 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[332] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__13_  ( .D(
        \iRF_stage/reg_bank/n471 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[333] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__14_  ( .D(
        \iRF_stage/reg_bank/n472 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[334] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__15_  ( .D(
        \iRF_stage/reg_bank/n473 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[335] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__16_  ( .D(
        \iRF_stage/reg_bank/n474 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[336] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__17_  ( .D(
        \iRF_stage/reg_bank/n475 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[337] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__18_  ( .D(
        \iRF_stage/reg_bank/n476 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[338] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__19_  ( .D(
        \iRF_stage/reg_bank/n477 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[339] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__20_  ( .D(
        \iRF_stage/reg_bank/n478 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[340] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__21_  ( .D(
        \iRF_stage/reg_bank/n479 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[341] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__22_  ( .D(
        \iRF_stage/reg_bank/n480 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[342] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__23_  ( .D(
        \iRF_stage/reg_bank/n481 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[343] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__24_  ( .D(
        \iRF_stage/reg_bank/n482 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[344] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__25_  ( .D(
        \iRF_stage/reg_bank/n483 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[345] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__26_  ( .D(
        \iRF_stage/reg_bank/n484 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[346] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__27_  ( .D(
        \iRF_stage/reg_bank/n485 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[347] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__28_  ( .D(
        \iRF_stage/reg_bank/n486 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[348] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__29_  ( .D(
        \iRF_stage/reg_bank/n487 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[349] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__30_  ( .D(
        \iRF_stage/reg_bank/n488 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[350] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_21__31_  ( .D(
        \iRF_stage/reg_bank/n489 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[351] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__0_  ( .D(
        \iRF_stage/reg_bank/n586 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[448] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__1_  ( .D(
        \iRF_stage/reg_bank/n587 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[449] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__2_  ( .D(
        \iRF_stage/reg_bank/n588 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[450] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__3_  ( .D(
        \iRF_stage/reg_bank/n589 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[451] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__4_  ( .D(
        \iRF_stage/reg_bank/n590 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[452] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__5_  ( .D(
        \iRF_stage/reg_bank/n591 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[453] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__6_  ( .D(
        \iRF_stage/reg_bank/n592 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[454] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__7_  ( .D(
        \iRF_stage/reg_bank/n593 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[455] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__8_  ( .D(
        \iRF_stage/reg_bank/n594 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[456] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__9_  ( .D(
        \iRF_stage/reg_bank/n595 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[457] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__10_  ( .D(
        \iRF_stage/reg_bank/n596 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[458] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__11_  ( .D(
        \iRF_stage/reg_bank/n597 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[459] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__12_  ( .D(
        \iRF_stage/reg_bank/n598 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[460] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__13_  ( .D(
        \iRF_stage/reg_bank/n599 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[461] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__14_  ( .D(
        \iRF_stage/reg_bank/n600 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[462] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__15_  ( .D(
        \iRF_stage/reg_bank/n601 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[463] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__16_  ( .D(
        \iRF_stage/reg_bank/n602 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[464] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__17_  ( .D(
        \iRF_stage/reg_bank/n603 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[465] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__18_  ( .D(
        \iRF_stage/reg_bank/n604 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[466] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__19_  ( .D(
        \iRF_stage/reg_bank/n605 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[467] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__20_  ( .D(
        \iRF_stage/reg_bank/n606 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[468] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__21_  ( .D(
        \iRF_stage/reg_bank/n607 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[469] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__22_  ( .D(
        \iRF_stage/reg_bank/n608 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[470] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__23_  ( .D(
        \iRF_stage/reg_bank/n609 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[471] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__24_  ( .D(
        \iRF_stage/reg_bank/n610 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[472] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__25_  ( .D(
        \iRF_stage/reg_bank/n611 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[473] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__26_  ( .D(
        \iRF_stage/reg_bank/n612 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[474] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__27_  ( .D(
        \iRF_stage/reg_bank/n613 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[475] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__28_  ( .D(
        \iRF_stage/reg_bank/n614 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[476] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__29_  ( .D(
        \iRF_stage/reg_bank/n615 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[477] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__30_  ( .D(
        \iRF_stage/reg_bank/n616 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[478] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_17__31_  ( .D(
        \iRF_stage/reg_bank/n617 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[479] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__0_  ( .D(
        \iRF_stage/reg_bank/n714 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[576] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__1_  ( .D(
        \iRF_stage/reg_bank/n715 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[577] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__2_  ( .D(
        \iRF_stage/reg_bank/n716 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[578] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__3_  ( .D(
        \iRF_stage/reg_bank/n717 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[579] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__4_  ( .D(
        \iRF_stage/reg_bank/n718 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[580] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__5_  ( .D(
        \iRF_stage/reg_bank/n719 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[581] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__6_  ( .D(
        \iRF_stage/reg_bank/n720 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[582] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__7_  ( .D(
        \iRF_stage/reg_bank/n721 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[583] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__8_  ( .D(
        \iRF_stage/reg_bank/n722 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[584] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__9_  ( .D(
        \iRF_stage/reg_bank/n723 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[585] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__10_  ( .D(
        \iRF_stage/reg_bank/n724 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[586] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__11_  ( .D(
        \iRF_stage/reg_bank/n725 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[587] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__12_  ( .D(
        \iRF_stage/reg_bank/n726 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[588] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__13_  ( .D(
        \iRF_stage/reg_bank/n727 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[589] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__14_  ( .D(
        \iRF_stage/reg_bank/n728 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[590] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__15_  ( .D(
        \iRF_stage/reg_bank/n729 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[591] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__16_  ( .D(
        \iRF_stage/reg_bank/n730 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[592] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__17_  ( .D(
        \iRF_stage/reg_bank/n731 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[593] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__18_  ( .D(
        \iRF_stage/reg_bank/n732 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[594] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__19_  ( .D(
        \iRF_stage/reg_bank/n733 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[595] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__20_  ( .D(
        \iRF_stage/reg_bank/n734 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[596] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__21_  ( .D(
        \iRF_stage/reg_bank/n735 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[597] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__22_  ( .D(
        \iRF_stage/reg_bank/n736 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[598] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__23_  ( .D(
        \iRF_stage/reg_bank/n737 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[599] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__24_  ( .D(
        \iRF_stage/reg_bank/n738 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[600] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__25_  ( .D(
        \iRF_stage/reg_bank/n739 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[601] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__26_  ( .D(
        \iRF_stage/reg_bank/n740 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[602] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__27_  ( .D(
        \iRF_stage/reg_bank/n741 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[603] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__28_  ( .D(
        \iRF_stage/reg_bank/n742 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[604] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__29_  ( .D(
        \iRF_stage/reg_bank/n743 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[605] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__30_  ( .D(
        \iRF_stage/reg_bank/n744 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[606] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_13__31_  ( .D(
        \iRF_stage/reg_bank/n745 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[607] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__0_  ( .D(
        \iRF_stage/reg_bank/n842 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[704] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__1_  ( .D(
        \iRF_stage/reg_bank/n843 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[705] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__2_  ( .D(
        \iRF_stage/reg_bank/n844 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[706] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__3_  ( .D(
        \iRF_stage/reg_bank/n845 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[707] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__4_  ( .D(
        \iRF_stage/reg_bank/n846 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[708] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__5_  ( .D(
        \iRF_stage/reg_bank/n847 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[709] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__6_  ( .D(
        \iRF_stage/reg_bank/n848 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[710] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__7_  ( .D(
        \iRF_stage/reg_bank/n849 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[711] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__8_  ( .D(
        \iRF_stage/reg_bank/n850 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[712] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__9_  ( .D(
        \iRF_stage/reg_bank/n851 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[713] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__10_  ( .D(
        \iRF_stage/reg_bank/n852 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[714] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__11_  ( .D(
        \iRF_stage/reg_bank/n853 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[715] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__12_  ( .D(
        \iRF_stage/reg_bank/n854 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[716] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__13_  ( .D(
        \iRF_stage/reg_bank/n855 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[717] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__14_  ( .D(
        \iRF_stage/reg_bank/n856 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[718] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__15_  ( .D(
        \iRF_stage/reg_bank/n857 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[719] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__16_  ( .D(
        \iRF_stage/reg_bank/n858 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[720] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__17_  ( .D(
        \iRF_stage/reg_bank/n859 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[721] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__18_  ( .D(
        \iRF_stage/reg_bank/n860 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[722] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__19_  ( .D(
        \iRF_stage/reg_bank/n861 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[723] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__20_  ( .D(
        \iRF_stage/reg_bank/n862 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[724] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__21_  ( .D(
        \iRF_stage/reg_bank/n863 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[725] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__22_  ( .D(
        \iRF_stage/reg_bank/n864 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[726] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__23_  ( .D(
        \iRF_stage/reg_bank/n865 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[727] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__24_  ( .D(
        \iRF_stage/reg_bank/n866 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[728] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__25_  ( .D(
        \iRF_stage/reg_bank/n867 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[729] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__26_  ( .D(
        \iRF_stage/reg_bank/n868 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[730] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__27_  ( .D(
        \iRF_stage/reg_bank/n869 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[731] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__28_  ( .D(
        \iRF_stage/reg_bank/n870 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[732] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__29_  ( .D(
        \iRF_stage/reg_bank/n871 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[733] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__30_  ( .D(
        \iRF_stage/reg_bank/n872 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[734] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_9__31_  ( .D(
        \iRF_stage/reg_bank/n873 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[735] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__0_  ( .D(
        \iRF_stage/reg_bank/n970 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[832] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__1_  ( .D(
        \iRF_stage/reg_bank/n971 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[833] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__2_  ( .D(
        \iRF_stage/reg_bank/n972 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[834] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__3_  ( .D(
        \iRF_stage/reg_bank/n973 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[835] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__4_  ( .D(
        \iRF_stage/reg_bank/n974 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[836] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__5_  ( .D(
        \iRF_stage/reg_bank/n975 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[837] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__6_  ( .D(
        \iRF_stage/reg_bank/n976 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[838] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__7_  ( .D(
        \iRF_stage/reg_bank/n977 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[839] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__8_  ( .D(
        \iRF_stage/reg_bank/n978 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[840] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__9_  ( .D(
        \iRF_stage/reg_bank/n979 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[841] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__10_  ( .D(
        \iRF_stage/reg_bank/n980 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[842] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__11_  ( .D(
        \iRF_stage/reg_bank/n981 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[843] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__12_  ( .D(
        \iRF_stage/reg_bank/n982 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[844] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__13_  ( .D(
        \iRF_stage/reg_bank/n983 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[845] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__14_  ( .D(
        \iRF_stage/reg_bank/n984 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[846] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__15_  ( .D(
        \iRF_stage/reg_bank/n985 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[847] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__16_  ( .D(
        \iRF_stage/reg_bank/n986 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[848] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__17_  ( .D(
        \iRF_stage/reg_bank/n987 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[849] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__18_  ( .D(
        \iRF_stage/reg_bank/n988 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[850] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__19_  ( .D(
        \iRF_stage/reg_bank/n989 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[851] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__20_  ( .D(
        \iRF_stage/reg_bank/n990 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[852] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__21_  ( .D(
        \iRF_stage/reg_bank/n991 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[853] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__22_  ( .D(
        \iRF_stage/reg_bank/n992 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[854] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__23_  ( .D(
        \iRF_stage/reg_bank/n993 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[855] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__24_  ( .D(
        \iRF_stage/reg_bank/n994 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[856] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__25_  ( .D(
        \iRF_stage/reg_bank/n995 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[857] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__26_  ( .D(
        \iRF_stage/reg_bank/n996 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[858] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__27_  ( .D(
        \iRF_stage/reg_bank/n997 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[859] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__28_  ( .D(
        \iRF_stage/reg_bank/n998 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[860] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__29_  ( .D(
        \iRF_stage/reg_bank/n999 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[861] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__30_  ( .D(
        \iRF_stage/reg_bank/n1000 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[862] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_5__31_  ( .D(
        \iRF_stage/reg_bank/n1001 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[863] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__0_  ( .D(
        \iRF_stage/reg_bank/n1098 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[960] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__1_  ( .D(
        \iRF_stage/reg_bank/n1099 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[961] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__2_  ( .D(
        \iRF_stage/reg_bank/n1100 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[962] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__3_  ( .D(
        \iRF_stage/reg_bank/n1101 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[963] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__4_  ( .D(
        \iRF_stage/reg_bank/n1102 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[964] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__5_  ( .D(
        \iRF_stage/reg_bank/n1103 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[965] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__6_  ( .D(
        \iRF_stage/reg_bank/n1104 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[966] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__7_  ( .D(
        \iRF_stage/reg_bank/n1105 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[967] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__8_  ( .D(
        \iRF_stage/reg_bank/n1106 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[968] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__9_  ( .D(
        \iRF_stage/reg_bank/n1107 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[969] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__10_  ( .D(
        \iRF_stage/reg_bank/n1108 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[970] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__11_  ( .D(
        \iRF_stage/reg_bank/n1109 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[971] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__12_  ( .D(
        \iRF_stage/reg_bank/n1110 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[972] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__13_  ( .D(
        \iRF_stage/reg_bank/n1111 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[973] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__14_  ( .D(
        \iRF_stage/reg_bank/n1112 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[974] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__15_  ( .D(
        \iRF_stage/reg_bank/n1113 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[975] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__16_  ( .D(
        \iRF_stage/reg_bank/n1114 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[976] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__17_  ( .D(
        \iRF_stage/reg_bank/n1115 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[977] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__18_  ( .D(
        \iRF_stage/reg_bank/n1116 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[978] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__19_  ( .D(
        \iRF_stage/reg_bank/n1117 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[979] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__20_  ( .D(
        \iRF_stage/reg_bank/n1118 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[980] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__21_  ( .D(
        \iRF_stage/reg_bank/n1119 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[981] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__22_  ( .D(
        \iRF_stage/reg_bank/n1120 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[982] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__23_  ( .D(
        \iRF_stage/reg_bank/n1121 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[983] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__24_  ( .D(
        \iRF_stage/reg_bank/n1122 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[984] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__25_  ( .D(
        \iRF_stage/reg_bank/n1123 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[985] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__26_  ( .D(
        \iRF_stage/reg_bank/n1124 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[986] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__27_  ( .D(
        \iRF_stage/reg_bank/n1125 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[987] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__28_  ( .D(
        \iRF_stage/reg_bank/n1126 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[988] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__29_  ( .D(
        \iRF_stage/reg_bank/n1127 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[989] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__30_  ( .D(
        \iRF_stage/reg_bank/n1128 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[990] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_1__31_  ( .D(
        \iRF_stage/reg_bank/n1129 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[991] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__0_  ( .D(
        \iRF_stage/reg_bank/n234 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[96] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__1_  ( .D(
        \iRF_stage/reg_bank/n235 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[97] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__2_  ( .D(
        \iRF_stage/reg_bank/n236 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[98] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__3_  ( .D(
        \iRF_stage/reg_bank/n237 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[99] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__4_  ( .D(
        \iRF_stage/reg_bank/n238 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[100] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__5_  ( .D(
        \iRF_stage/reg_bank/n239 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[101] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__6_  ( .D(
        \iRF_stage/reg_bank/n240 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[102] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__7_  ( .D(
        \iRF_stage/reg_bank/n241 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[103] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__8_  ( .D(
        \iRF_stage/reg_bank/n242 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[104] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__9_  ( .D(
        \iRF_stage/reg_bank/n243 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[105] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__10_  ( .D(
        \iRF_stage/reg_bank/n244 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[106] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__11_  ( .D(
        \iRF_stage/reg_bank/n245 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[107] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__12_  ( .D(
        \iRF_stage/reg_bank/n246 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[108] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__13_  ( .D(
        \iRF_stage/reg_bank/n247 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[109] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__14_  ( .D(
        \iRF_stage/reg_bank/n248 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[110] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__15_  ( .D(
        \iRF_stage/reg_bank/n249 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[111] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__16_  ( .D(
        \iRF_stage/reg_bank/n250 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[112] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__17_  ( .D(
        \iRF_stage/reg_bank/n251 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[113] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__18_  ( .D(
        \iRF_stage/reg_bank/n252 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[114] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__19_  ( .D(
        \iRF_stage/reg_bank/n253 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[115] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__20_  ( .D(
        \iRF_stage/reg_bank/n254 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[116] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__21_  ( .D(
        \iRF_stage/reg_bank/n255 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[117] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__22_  ( .D(
        \iRF_stage/reg_bank/n256 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[118] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__23_  ( .D(
        \iRF_stage/reg_bank/n257 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[119] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__24_  ( .D(
        \iRF_stage/reg_bank/n258 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[120] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__25_  ( .D(
        \iRF_stage/reg_bank/n259 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[121] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__26_  ( .D(
        \iRF_stage/reg_bank/n260 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[122] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__27_  ( .D(
        \iRF_stage/reg_bank/n261 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[123] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__28_  ( .D(
        \iRF_stage/reg_bank/n262 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[124] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__29_  ( .D(
        \iRF_stage/reg_bank/n263 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[125] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__30_  ( .D(
        \iRF_stage/reg_bank/n264 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[126] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_28__31_  ( .D(
        \iRF_stage/reg_bank/n265 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[127] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__0_  ( .D(
        \iRF_stage/reg_bank/n362 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[224] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__1_  ( .D(
        \iRF_stage/reg_bank/n363 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[225] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__2_  ( .D(
        \iRF_stage/reg_bank/n364 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[226] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__3_  ( .D(
        \iRF_stage/reg_bank/n365 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[227] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__4_  ( .D(
        \iRF_stage/reg_bank/n366 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[228] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__5_  ( .D(
        \iRF_stage/reg_bank/n367 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[229] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__6_  ( .D(
        \iRF_stage/reg_bank/n368 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[230] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__7_  ( .D(
        \iRF_stage/reg_bank/n369 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[231] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__8_  ( .D(
        \iRF_stage/reg_bank/n370 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[232] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__9_  ( .D(
        \iRF_stage/reg_bank/n371 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[233] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__10_  ( .D(
        \iRF_stage/reg_bank/n372 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[234] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__11_  ( .D(
        \iRF_stage/reg_bank/n373 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[235] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__12_  ( .D(
        \iRF_stage/reg_bank/n374 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[236] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__13_  ( .D(
        \iRF_stage/reg_bank/n375 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[237] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__14_  ( .D(
        \iRF_stage/reg_bank/n376 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[238] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__15_  ( .D(
        \iRF_stage/reg_bank/n377 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[239] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__16_  ( .D(
        \iRF_stage/reg_bank/n378 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[240] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__17_  ( .D(
        \iRF_stage/reg_bank/n379 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[241] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__18_  ( .D(
        \iRF_stage/reg_bank/n380 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[242] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__19_  ( .D(
        \iRF_stage/reg_bank/n381 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[243] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__20_  ( .D(
        \iRF_stage/reg_bank/n382 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[244] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__21_  ( .D(
        \iRF_stage/reg_bank/n383 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[245] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__22_  ( .D(
        \iRF_stage/reg_bank/n384 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[246] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__23_  ( .D(
        \iRF_stage/reg_bank/n385 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[247] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__24_  ( .D(
        \iRF_stage/reg_bank/n386 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[248] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__25_  ( .D(
        \iRF_stage/reg_bank/n387 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[249] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__26_  ( .D(
        \iRF_stage/reg_bank/n388 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[250] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__27_  ( .D(
        \iRF_stage/reg_bank/n389 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[251] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__28_  ( .D(
        \iRF_stage/reg_bank/n390 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[252] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__29_  ( .D(
        \iRF_stage/reg_bank/n391 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[253] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__30_  ( .D(
        \iRF_stage/reg_bank/n392 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[254] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_24__31_  ( .D(
        \iRF_stage/reg_bank/n393 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[255] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__0_  ( .D(
        \iRF_stage/reg_bank/n490 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[352] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__1_  ( .D(
        \iRF_stage/reg_bank/n491 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[353] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__2_  ( .D(
        \iRF_stage/reg_bank/n492 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[354] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__3_  ( .D(
        \iRF_stage/reg_bank/n493 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[355] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__4_  ( .D(
        \iRF_stage/reg_bank/n494 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[356] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__5_  ( .D(
        \iRF_stage/reg_bank/n495 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[357] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__6_  ( .D(
        \iRF_stage/reg_bank/n496 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[358] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__7_  ( .D(
        \iRF_stage/reg_bank/n497 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[359] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__8_  ( .D(
        \iRF_stage/reg_bank/n498 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[360] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__9_  ( .D(
        \iRF_stage/reg_bank/n499 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[361] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__10_  ( .D(
        \iRF_stage/reg_bank/n500 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[362] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__11_  ( .D(
        \iRF_stage/reg_bank/n501 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[363] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__12_  ( .D(
        \iRF_stage/reg_bank/n502 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[364] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__13_  ( .D(
        \iRF_stage/reg_bank/n503 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[365] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__14_  ( .D(
        \iRF_stage/reg_bank/n504 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[366] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__15_  ( .D(
        \iRF_stage/reg_bank/n505 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[367] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__16_  ( .D(
        \iRF_stage/reg_bank/n506 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[368] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__17_  ( .D(
        \iRF_stage/reg_bank/n507 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[369] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__18_  ( .D(
        \iRF_stage/reg_bank/n508 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[370] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__19_  ( .D(
        \iRF_stage/reg_bank/n509 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[371] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__20_  ( .D(
        \iRF_stage/reg_bank/n510 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[372] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__21_  ( .D(
        \iRF_stage/reg_bank/n511 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[373] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__22_  ( .D(
        \iRF_stage/reg_bank/n512 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[374] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__23_  ( .D(
        \iRF_stage/reg_bank/n513 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[375] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__24_  ( .D(
        \iRF_stage/reg_bank/n514 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[376] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__25_  ( .D(
        \iRF_stage/reg_bank/n515 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[377] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__26_  ( .D(
        \iRF_stage/reg_bank/n516 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[378] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__27_  ( .D(
        \iRF_stage/reg_bank/n517 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[379] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__28_  ( .D(
        \iRF_stage/reg_bank/n518 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[380] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__29_  ( .D(
        \iRF_stage/reg_bank/n519 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[381] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__30_  ( .D(
        \iRF_stage/reg_bank/n520 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[382] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_20__31_  ( .D(
        \iRF_stage/reg_bank/n521 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[383] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__0_  ( .D(
        \iRF_stage/reg_bank/n618 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[480] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__1_  ( .D(
        \iRF_stage/reg_bank/n619 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[481] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__2_  ( .D(
        \iRF_stage/reg_bank/n620 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[482] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__3_  ( .D(
        \iRF_stage/reg_bank/n621 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[483] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__4_  ( .D(
        \iRF_stage/reg_bank/n622 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[484] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__5_  ( .D(
        \iRF_stage/reg_bank/n623 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[485] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__6_  ( .D(
        \iRF_stage/reg_bank/n624 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[486] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__7_  ( .D(
        \iRF_stage/reg_bank/n625 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[487] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__8_  ( .D(
        \iRF_stage/reg_bank/n626 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[488] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__9_  ( .D(
        \iRF_stage/reg_bank/n627 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[489] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__10_  ( .D(
        \iRF_stage/reg_bank/n628 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[490] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__11_  ( .D(
        \iRF_stage/reg_bank/n629 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[491] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__12_  ( .D(
        \iRF_stage/reg_bank/n630 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[492] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__13_  ( .D(
        \iRF_stage/reg_bank/n631 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[493] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__14_  ( .D(
        \iRF_stage/reg_bank/n632 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[494] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__15_  ( .D(
        \iRF_stage/reg_bank/n633 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[495] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__16_  ( .D(
        \iRF_stage/reg_bank/n634 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[496] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__17_  ( .D(
        \iRF_stage/reg_bank/n635 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[497] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__18_  ( .D(
        \iRF_stage/reg_bank/n636 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[498] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__19_  ( .D(
        \iRF_stage/reg_bank/n637 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[499] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__20_  ( .D(
        \iRF_stage/reg_bank/n638 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[500] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__21_  ( .D(
        \iRF_stage/reg_bank/n639 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[501] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__22_  ( .D(
        \iRF_stage/reg_bank/n640 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[502] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__23_  ( .D(
        \iRF_stage/reg_bank/n641 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[503] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__24_  ( .D(
        \iRF_stage/reg_bank/n642 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[504] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__25_  ( .D(
        \iRF_stage/reg_bank/n643 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[505] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__26_  ( .D(
        \iRF_stage/reg_bank/n644 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[506] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__27_  ( .D(
        \iRF_stage/reg_bank/n645 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[507] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__28_  ( .D(
        \iRF_stage/reg_bank/n646 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[508] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__29_  ( .D(
        \iRF_stage/reg_bank/n647 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[509] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__30_  ( .D(
        \iRF_stage/reg_bank/n648 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[510] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_16__31_  ( .D(
        \iRF_stage/reg_bank/n649 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[511] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__0_  ( .D(
        \iRF_stage/reg_bank/n746 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[608] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__1_  ( .D(
        \iRF_stage/reg_bank/n747 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[609] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__2_  ( .D(
        \iRF_stage/reg_bank/n748 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[610] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__3_  ( .D(
        \iRF_stage/reg_bank/n749 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[611] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__4_  ( .D(
        \iRF_stage/reg_bank/n750 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[612] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__5_  ( .D(
        \iRF_stage/reg_bank/n751 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[613] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__6_  ( .D(
        \iRF_stage/reg_bank/n752 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[614] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__7_  ( .D(
        \iRF_stage/reg_bank/n753 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[615] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__8_  ( .D(
        \iRF_stage/reg_bank/n754 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[616] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__9_  ( .D(
        \iRF_stage/reg_bank/n755 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[617] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__10_  ( .D(
        \iRF_stage/reg_bank/n756 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[618] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__11_  ( .D(
        \iRF_stage/reg_bank/n757 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[619] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__12_  ( .D(
        \iRF_stage/reg_bank/n758 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[620] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__13_  ( .D(
        \iRF_stage/reg_bank/n759 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[621] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__14_  ( .D(
        \iRF_stage/reg_bank/n760 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[622] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__15_  ( .D(
        \iRF_stage/reg_bank/n761 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[623] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__16_  ( .D(
        \iRF_stage/reg_bank/n762 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[624] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__17_  ( .D(
        \iRF_stage/reg_bank/n763 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[625] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__18_  ( .D(
        \iRF_stage/reg_bank/n764 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[626] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__19_  ( .D(
        \iRF_stage/reg_bank/n765 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[627] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__20_  ( .D(
        \iRF_stage/reg_bank/n766 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[628] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__21_  ( .D(
        \iRF_stage/reg_bank/n767 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[629] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__22_  ( .D(
        \iRF_stage/reg_bank/n768 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[630] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__23_  ( .D(
        \iRF_stage/reg_bank/n769 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[631] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__24_  ( .D(
        \iRF_stage/reg_bank/n770 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[632] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__25_  ( .D(
        \iRF_stage/reg_bank/n771 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[633] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__26_  ( .D(
        \iRF_stage/reg_bank/n772 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[634] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__27_  ( .D(
        \iRF_stage/reg_bank/n773 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[635] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__28_  ( .D(
        \iRF_stage/reg_bank/n774 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[636] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__29_  ( .D(
        \iRF_stage/reg_bank/n775 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[637] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__30_  ( .D(
        \iRF_stage/reg_bank/n776 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[638] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_12__31_  ( .D(
        \iRF_stage/reg_bank/n777 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[639] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__0_  ( .D(
        \iRF_stage/reg_bank/n874 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[736] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__1_  ( .D(
        \iRF_stage/reg_bank/n875 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[737] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__2_  ( .D(
        \iRF_stage/reg_bank/n876 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[738] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__3_  ( .D(
        \iRF_stage/reg_bank/n877 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[739] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__4_  ( .D(
        \iRF_stage/reg_bank/n878 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[740] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__5_  ( .D(
        \iRF_stage/reg_bank/n879 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[741] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__6_  ( .D(
        \iRF_stage/reg_bank/n880 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[742] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__7_  ( .D(
        \iRF_stage/reg_bank/n881 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[743] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__8_  ( .D(
        \iRF_stage/reg_bank/n882 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[744] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__9_  ( .D(
        \iRF_stage/reg_bank/n883 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[745] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__10_  ( .D(
        \iRF_stage/reg_bank/n884 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[746] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__11_  ( .D(
        \iRF_stage/reg_bank/n885 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[747] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__12_  ( .D(
        \iRF_stage/reg_bank/n886 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[748] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__13_  ( .D(
        \iRF_stage/reg_bank/n887 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[749] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__14_  ( .D(
        \iRF_stage/reg_bank/n888 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[750] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__15_  ( .D(
        \iRF_stage/reg_bank/n889 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[751] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__16_  ( .D(
        \iRF_stage/reg_bank/n890 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[752] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__17_  ( .D(
        \iRF_stage/reg_bank/n891 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[753] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__18_  ( .D(
        \iRF_stage/reg_bank/n892 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[754] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__19_  ( .D(
        \iRF_stage/reg_bank/n893 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[755] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__20_  ( .D(
        \iRF_stage/reg_bank/n894 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[756] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__21_  ( .D(
        \iRF_stage/reg_bank/n895 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[757] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__22_  ( .D(
        \iRF_stage/reg_bank/n896 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[758] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__23_  ( .D(
        \iRF_stage/reg_bank/n897 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[759] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__24_  ( .D(
        \iRF_stage/reg_bank/n898 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[760] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__25_  ( .D(
        \iRF_stage/reg_bank/n899 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[761] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__26_  ( .D(
        \iRF_stage/reg_bank/n900 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[762] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__27_  ( .D(
        \iRF_stage/reg_bank/n901 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[763] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__28_  ( .D(
        \iRF_stage/reg_bank/n902 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[764] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__29_  ( .D(
        \iRF_stage/reg_bank/n903 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[765] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__30_  ( .D(
        \iRF_stage/reg_bank/n904 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[766] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_8__31_  ( .D(
        \iRF_stage/reg_bank/n905 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[767] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__0_  ( .D(
        \iRF_stage/reg_bank/n1002 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[864] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__1_  ( .D(
        \iRF_stage/reg_bank/n1003 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[865] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__2_  ( .D(
        \iRF_stage/reg_bank/n1004 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[866] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__3_  ( .D(
        \iRF_stage/reg_bank/n1005 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[867] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__4_  ( .D(
        \iRF_stage/reg_bank/n1006 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[868] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__5_  ( .D(
        \iRF_stage/reg_bank/n1007 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[869] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__6_  ( .D(
        \iRF_stage/reg_bank/n1008 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[870] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__7_  ( .D(
        \iRF_stage/reg_bank/n1009 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[871] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__8_  ( .D(
        \iRF_stage/reg_bank/n1010 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[872] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__9_  ( .D(
        \iRF_stage/reg_bank/n1011 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[873] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__10_  ( .D(
        \iRF_stage/reg_bank/n1012 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[874] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__11_  ( .D(
        \iRF_stage/reg_bank/n1013 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[875] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__12_  ( .D(
        \iRF_stage/reg_bank/n1014 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[876] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__13_  ( .D(
        \iRF_stage/reg_bank/n1015 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[877] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__14_  ( .D(
        \iRF_stage/reg_bank/n1016 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[878] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__15_  ( .D(
        \iRF_stage/reg_bank/n1017 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[879] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__16_  ( .D(
        \iRF_stage/reg_bank/n1018 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[880] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__17_  ( .D(
        \iRF_stage/reg_bank/n1019 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[881] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__18_  ( .D(
        \iRF_stage/reg_bank/n1020 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[882] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__19_  ( .D(
        \iRF_stage/reg_bank/n1021 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[883] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__20_  ( .D(
        \iRF_stage/reg_bank/n1022 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[884] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__21_  ( .D(
        \iRF_stage/reg_bank/n1023 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[885] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__22_  ( .D(
        \iRF_stage/reg_bank/n1024 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[886] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__23_  ( .D(
        \iRF_stage/reg_bank/n1025 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[887] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__24_  ( .D(
        \iRF_stage/reg_bank/n1026 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[888] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__25_  ( .D(
        \iRF_stage/reg_bank/n1027 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[889] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__26_  ( .D(
        \iRF_stage/reg_bank/n1028 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[890] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__27_  ( .D(
        \iRF_stage/reg_bank/n1029 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[891] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__28_  ( .D(
        \iRF_stage/reg_bank/n1030 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[892] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__29_  ( .D(
        \iRF_stage/reg_bank/n1031 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[893] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__30_  ( .D(
        \iRF_stage/reg_bank/n1032 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[894] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_4__31_  ( .D(
        \iRF_stage/reg_bank/n1033 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[895] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__0_  ( .D(
        \iRF_stage/reg_bank/n1130 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[992] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__1_  ( .D(
        \iRF_stage/reg_bank/n1131 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[993] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__2_  ( .D(
        \iRF_stage/reg_bank/n1132 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[994] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__3_  ( .D(
        \iRF_stage/reg_bank/n1133 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[995] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__4_  ( .D(
        \iRF_stage/reg_bank/n1134 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[996] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__5_  ( .D(
        \iRF_stage/reg_bank/n1135 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[997] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__6_  ( .D(
        \iRF_stage/reg_bank/n1136 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[998] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__7_  ( .D(
        \iRF_stage/reg_bank/n1137 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[999] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__8_  ( .D(
        \iRF_stage/reg_bank/n1138 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1000] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__9_  ( .D(
        \iRF_stage/reg_bank/n1139 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1001] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__10_  ( .D(
        \iRF_stage/reg_bank/n1140 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1002] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__11_  ( .D(
        \iRF_stage/reg_bank/n1141 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1003] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__12_  ( .D(
        \iRF_stage/reg_bank/n1142 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1004] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__13_  ( .D(
        \iRF_stage/reg_bank/n1143 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1005] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__14_  ( .D(
        \iRF_stage/reg_bank/n1144 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1006] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__15_  ( .D(
        \iRF_stage/reg_bank/n1145 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1007] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__16_  ( .D(
        \iRF_stage/reg_bank/n1146 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1008] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__17_  ( .D(
        \iRF_stage/reg_bank/n1147 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1009] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__18_  ( .D(
        \iRF_stage/reg_bank/n1148 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1010] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__19_  ( .D(
        \iRF_stage/reg_bank/n1149 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1011] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__20_  ( .D(
        \iRF_stage/reg_bank/n1150 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1012] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__21_  ( .D(
        \iRF_stage/reg_bank/n1151 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1013] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__22_  ( .D(
        \iRF_stage/reg_bank/n1152 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1014] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__23_  ( .D(
        \iRF_stage/reg_bank/n1153 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1015] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__24_  ( .D(
        \iRF_stage/reg_bank/n1154 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1016] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__25_  ( .D(
        \iRF_stage/reg_bank/n1155 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1017] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__26_  ( .D(
        \iRF_stage/reg_bank/n1156 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1018] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__27_  ( .D(
        \iRF_stage/reg_bank/n1157 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1019] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__28_  ( .D(
        \iRF_stage/reg_bank/n1158 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1020] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__29_  ( .D(
        \iRF_stage/reg_bank/n1159 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1021] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__30_  ( .D(
        \iRF_stage/reg_bank/n1160 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1022] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_0__31_  ( .D(
        \iRF_stage/reg_bank/n1161 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1023] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__0_  ( .D(
        \iRF_stage/reg_bank/n138 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[0] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__1_  ( .D(
        \iRF_stage/reg_bank/n139 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[1] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__2_  ( .D(
        \iRF_stage/reg_bank/n140 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[2] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__3_  ( .D(
        \iRF_stage/reg_bank/n141 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[3] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__4_  ( .D(
        \iRF_stage/reg_bank/n142 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[4] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__5_  ( .D(
        \iRF_stage/reg_bank/n143 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[5] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__6_  ( .D(
        \iRF_stage/reg_bank/n144 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[6] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__7_  ( .D(
        \iRF_stage/reg_bank/n145 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[7] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__8_  ( .D(
        \iRF_stage/reg_bank/n146 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[8] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__9_  ( .D(
        \iRF_stage/reg_bank/n147 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[9] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__10_  ( .D(
        \iRF_stage/reg_bank/n148 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[10] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__11_  ( .D(
        \iRF_stage/reg_bank/n149 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[11] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__12_  ( .D(
        \iRF_stage/reg_bank/n150 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[12] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__13_  ( .D(
        \iRF_stage/reg_bank/n151 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[13] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__14_  ( .D(
        \iRF_stage/reg_bank/n152 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[14] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__15_  ( .D(
        \iRF_stage/reg_bank/n153 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[15] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__16_  ( .D(
        \iRF_stage/reg_bank/n154 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[16] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__17_  ( .D(
        \iRF_stage/reg_bank/n155 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[17] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__18_  ( .D(
        \iRF_stage/reg_bank/n156 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[18] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__19_  ( .D(
        \iRF_stage/reg_bank/n157 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[19] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__20_  ( .D(
        \iRF_stage/reg_bank/n158 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[20] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__21_  ( .D(
        \iRF_stage/reg_bank/n159 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[21] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__22_  ( .D(
        \iRF_stage/reg_bank/n160 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[22] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__23_  ( .D(
        \iRF_stage/reg_bank/n161 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[23] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__24_  ( .D(
        \iRF_stage/reg_bank/n162 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[24] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__25_  ( .D(
        \iRF_stage/reg_bank/n163 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[25] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__26_  ( .D(
        \iRF_stage/reg_bank/n164 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[26] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__27_  ( .D(
        \iRF_stage/reg_bank/n165 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[27] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__28_  ( .D(
        \iRF_stage/reg_bank/n166 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[28] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__29_  ( .D(
        \iRF_stage/reg_bank/n167 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[29] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__30_  ( .D(
        \iRF_stage/reg_bank/n168 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[30] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_31__31_  ( .D(
        \iRF_stage/reg_bank/n169 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[31] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__0_  ( .D(
        \iRF_stage/reg_bank/n266 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[128] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__1_  ( .D(
        \iRF_stage/reg_bank/n267 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[129] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__2_  ( .D(
        \iRF_stage/reg_bank/n268 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[130] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__3_  ( .D(
        \iRF_stage/reg_bank/n269 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[131] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__4_  ( .D(
        \iRF_stage/reg_bank/n270 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[132] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__5_  ( .D(
        \iRF_stage/reg_bank/n271 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[133] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__6_  ( .D(
        \iRF_stage/reg_bank/n272 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[134] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__7_  ( .D(
        \iRF_stage/reg_bank/n273 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[135] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__8_  ( .D(
        \iRF_stage/reg_bank/n274 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[136] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__9_  ( .D(
        \iRF_stage/reg_bank/n275 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[137] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__10_  ( .D(
        \iRF_stage/reg_bank/n276 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[138] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__11_  ( .D(
        \iRF_stage/reg_bank/n277 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[139] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__12_  ( .D(
        \iRF_stage/reg_bank/n278 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[140] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__13_  ( .D(
        \iRF_stage/reg_bank/n279 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[141] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__14_  ( .D(
        \iRF_stage/reg_bank/n280 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[142] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__15_  ( .D(
        \iRF_stage/reg_bank/n281 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[143] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__16_  ( .D(
        \iRF_stage/reg_bank/n282 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[144] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__17_  ( .D(
        \iRF_stage/reg_bank/n283 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[145] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__18_  ( .D(
        \iRF_stage/reg_bank/n284 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[146] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__19_  ( .D(
        \iRF_stage/reg_bank/n285 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[147] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__20_  ( .D(
        \iRF_stage/reg_bank/n286 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[148] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__21_  ( .D(
        \iRF_stage/reg_bank/n287 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[149] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__22_  ( .D(
        \iRF_stage/reg_bank/n288 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[150] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__23_  ( .D(
        \iRF_stage/reg_bank/n289 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[151] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__24_  ( .D(
        \iRF_stage/reg_bank/n290 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[152] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__25_  ( .D(
        \iRF_stage/reg_bank/n291 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[153] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__26_  ( .D(
        \iRF_stage/reg_bank/n292 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[154] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__27_  ( .D(
        \iRF_stage/reg_bank/n293 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[155] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__28_  ( .D(
        \iRF_stage/reg_bank/n294 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[156] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__29_  ( .D(
        \iRF_stage/reg_bank/n295 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[157] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__30_  ( .D(
        \iRF_stage/reg_bank/n296 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[158] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_27__31_  ( .D(
        \iRF_stage/reg_bank/n297 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[159] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__0_  ( .D(
        \iRF_stage/reg_bank/n394 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[256] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__1_  ( .D(
        \iRF_stage/reg_bank/n395 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[257] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__2_  ( .D(
        \iRF_stage/reg_bank/n396 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[258] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__3_  ( .D(
        \iRF_stage/reg_bank/n397 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[259] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__4_  ( .D(
        \iRF_stage/reg_bank/n398 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[260] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__5_  ( .D(
        \iRF_stage/reg_bank/n399 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[261] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__6_  ( .D(
        \iRF_stage/reg_bank/n400 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[262] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__7_  ( .D(
        \iRF_stage/reg_bank/n401 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[263] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__8_  ( .D(
        \iRF_stage/reg_bank/n402 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[264] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__9_  ( .D(
        \iRF_stage/reg_bank/n403 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[265] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__10_  ( .D(
        \iRF_stage/reg_bank/n404 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[266] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__11_  ( .D(
        \iRF_stage/reg_bank/n405 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[267] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__12_  ( .D(
        \iRF_stage/reg_bank/n406 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[268] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__13_  ( .D(
        \iRF_stage/reg_bank/n407 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[269] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__14_  ( .D(
        \iRF_stage/reg_bank/n408 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[270] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__15_  ( .D(
        \iRF_stage/reg_bank/n409 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[271] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__16_  ( .D(
        \iRF_stage/reg_bank/n410 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[272] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__17_  ( .D(
        \iRF_stage/reg_bank/n411 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[273] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__18_  ( .D(
        \iRF_stage/reg_bank/n412 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[274] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__19_  ( .D(
        \iRF_stage/reg_bank/n413 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[275] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__20_  ( .D(
        \iRF_stage/reg_bank/n414 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[276] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__21_  ( .D(
        \iRF_stage/reg_bank/n415 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[277] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__22_  ( .D(
        \iRF_stage/reg_bank/n416 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[278] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__23_  ( .D(
        \iRF_stage/reg_bank/n417 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[279] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__24_  ( .D(
        \iRF_stage/reg_bank/n418 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[280] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__25_  ( .D(
        \iRF_stage/reg_bank/n419 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[281] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__26_  ( .D(
        \iRF_stage/reg_bank/n420 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[282] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__27_  ( .D(
        \iRF_stage/reg_bank/n421 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[283] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__28_  ( .D(
        \iRF_stage/reg_bank/n422 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[284] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__29_  ( .D(
        \iRF_stage/reg_bank/n423 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[285] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__30_  ( .D(
        \iRF_stage/reg_bank/n424 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[286] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_23__31_  ( .D(
        \iRF_stage/reg_bank/n425 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[287] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__0_  ( .D(
        \iRF_stage/reg_bank/n522 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[384] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__1_  ( .D(
        \iRF_stage/reg_bank/n523 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[385] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__2_  ( .D(
        \iRF_stage/reg_bank/n524 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[386] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__3_  ( .D(
        \iRF_stage/reg_bank/n525 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[387] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__4_  ( .D(
        \iRF_stage/reg_bank/n526 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[388] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__5_  ( .D(
        \iRF_stage/reg_bank/n527 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[389] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__6_  ( .D(
        \iRF_stage/reg_bank/n528 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[390] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__7_  ( .D(
        \iRF_stage/reg_bank/n529 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[391] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__8_  ( .D(
        \iRF_stage/reg_bank/n530 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[392] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__9_  ( .D(
        \iRF_stage/reg_bank/n531 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[393] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__10_  ( .D(
        \iRF_stage/reg_bank/n532 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[394] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__11_  ( .D(
        \iRF_stage/reg_bank/n533 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[395] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__12_  ( .D(
        \iRF_stage/reg_bank/n534 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[396] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__13_  ( .D(
        \iRF_stage/reg_bank/n535 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[397] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__14_  ( .D(
        \iRF_stage/reg_bank/n536 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[398] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__15_  ( .D(
        \iRF_stage/reg_bank/n537 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[399] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__16_  ( .D(
        \iRF_stage/reg_bank/n538 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[400] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__17_  ( .D(
        \iRF_stage/reg_bank/n539 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[401] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__18_  ( .D(
        \iRF_stage/reg_bank/n540 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[402] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__19_  ( .D(
        \iRF_stage/reg_bank/n541 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[403] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__20_  ( .D(
        \iRF_stage/reg_bank/n542 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[404] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__21_  ( .D(
        \iRF_stage/reg_bank/n543 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[405] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__22_  ( .D(
        \iRF_stage/reg_bank/n544 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[406] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__23_  ( .D(
        \iRF_stage/reg_bank/n545 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[407] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__24_  ( .D(
        \iRF_stage/reg_bank/n546 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[408] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__25_  ( .D(
        \iRF_stage/reg_bank/n547 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[409] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__26_  ( .D(
        \iRF_stage/reg_bank/n548 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[410] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__27_  ( .D(
        \iRF_stage/reg_bank/n549 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[411] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__28_  ( .D(
        \iRF_stage/reg_bank/n550 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[412] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__29_  ( .D(
        \iRF_stage/reg_bank/n551 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[413] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__30_  ( .D(
        \iRF_stage/reg_bank/n552 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[414] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_19__31_  ( .D(
        \iRF_stage/reg_bank/n553 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[415] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__0_  ( .D(
        \iRF_stage/reg_bank/n650 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[512] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__1_  ( .D(
        \iRF_stage/reg_bank/n651 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[513] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__2_  ( .D(
        \iRF_stage/reg_bank/n652 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[514] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__3_  ( .D(
        \iRF_stage/reg_bank/n653 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[515] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__4_  ( .D(
        \iRF_stage/reg_bank/n654 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[516] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__5_  ( .D(
        \iRF_stage/reg_bank/n655 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[517] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__6_  ( .D(
        \iRF_stage/reg_bank/n656 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[518] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__7_  ( .D(
        \iRF_stage/reg_bank/n657 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[519] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__8_  ( .D(
        \iRF_stage/reg_bank/n658 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[520] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__9_  ( .D(
        \iRF_stage/reg_bank/n659 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[521] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__10_  ( .D(
        \iRF_stage/reg_bank/n660 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[522] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__11_  ( .D(
        \iRF_stage/reg_bank/n661 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[523] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__12_  ( .D(
        \iRF_stage/reg_bank/n662 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[524] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__13_  ( .D(
        \iRF_stage/reg_bank/n663 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[525] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__14_  ( .D(
        \iRF_stage/reg_bank/n664 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[526] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__15_  ( .D(
        \iRF_stage/reg_bank/n665 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[527] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__16_  ( .D(
        \iRF_stage/reg_bank/n666 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[528] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__17_  ( .D(
        \iRF_stage/reg_bank/n667 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[529] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__18_  ( .D(
        \iRF_stage/reg_bank/n668 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[530] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__19_  ( .D(
        \iRF_stage/reg_bank/n669 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[531] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__20_  ( .D(
        \iRF_stage/reg_bank/n670 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[532] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__21_  ( .D(
        \iRF_stage/reg_bank/n671 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[533] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__22_  ( .D(
        \iRF_stage/reg_bank/n672 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[534] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__23_  ( .D(
        \iRF_stage/reg_bank/n673 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[535] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__24_  ( .D(
        \iRF_stage/reg_bank/n674 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[536] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__25_  ( .D(
        \iRF_stage/reg_bank/n675 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[537] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__26_  ( .D(
        \iRF_stage/reg_bank/n676 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[538] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__27_  ( .D(
        \iRF_stage/reg_bank/n677 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[539] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__28_  ( .D(
        \iRF_stage/reg_bank/n678 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[540] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__29_  ( .D(
        \iRF_stage/reg_bank/n679 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[541] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__30_  ( .D(
        \iRF_stage/reg_bank/n680 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[542] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_15__31_  ( .D(
        \iRF_stage/reg_bank/n681 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[543] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__0_  ( .D(
        \iRF_stage/reg_bank/n778 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[640] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__1_  ( .D(
        \iRF_stage/reg_bank/n779 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[641] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__2_  ( .D(
        \iRF_stage/reg_bank/n780 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[642] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__3_  ( .D(
        \iRF_stage/reg_bank/n781 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[643] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__4_  ( .D(
        \iRF_stage/reg_bank/n782 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[644] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__5_  ( .D(
        \iRF_stage/reg_bank/n783 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[645] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__6_  ( .D(
        \iRF_stage/reg_bank/n784 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[646] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__7_  ( .D(
        \iRF_stage/reg_bank/n785 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[647] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__8_  ( .D(
        \iRF_stage/reg_bank/n786 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[648] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__9_  ( .D(
        \iRF_stage/reg_bank/n787 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[649] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__10_  ( .D(
        \iRF_stage/reg_bank/n788 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[650] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__11_  ( .D(
        \iRF_stage/reg_bank/n789 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[651] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__12_  ( .D(
        \iRF_stage/reg_bank/n790 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[652] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__13_  ( .D(
        \iRF_stage/reg_bank/n791 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[653] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__14_  ( .D(
        \iRF_stage/reg_bank/n792 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[654] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__15_  ( .D(
        \iRF_stage/reg_bank/n793 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[655] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__16_  ( .D(
        \iRF_stage/reg_bank/n794 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[656] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__17_  ( .D(
        \iRF_stage/reg_bank/n795 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[657] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__18_  ( .D(
        \iRF_stage/reg_bank/n796 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[658] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__19_  ( .D(
        \iRF_stage/reg_bank/n797 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[659] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__20_  ( .D(
        \iRF_stage/reg_bank/n798 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[660] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__21_  ( .D(
        \iRF_stage/reg_bank/n799 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[661] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__22_  ( .D(
        \iRF_stage/reg_bank/n800 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[662] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__23_  ( .D(
        \iRF_stage/reg_bank/n801 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[663] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__24_  ( .D(
        \iRF_stage/reg_bank/n802 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[664] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__25_  ( .D(
        \iRF_stage/reg_bank/n803 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[665] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__26_  ( .D(
        \iRF_stage/reg_bank/n804 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[666] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__27_  ( .D(
        \iRF_stage/reg_bank/n805 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[667] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__28_  ( .D(
        \iRF_stage/reg_bank/n806 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[668] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__29_  ( .D(
        \iRF_stage/reg_bank/n807 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[669] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__30_  ( .D(
        \iRF_stage/reg_bank/n808 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[670] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_11__31_  ( .D(
        \iRF_stage/reg_bank/n809 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[671] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__0_  ( .D(
        \iRF_stage/reg_bank/n906 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[768] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__1_  ( .D(
        \iRF_stage/reg_bank/n907 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[769] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__2_  ( .D(
        \iRF_stage/reg_bank/n908 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[770] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__3_  ( .D(
        \iRF_stage/reg_bank/n909 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[771] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__4_  ( .D(
        \iRF_stage/reg_bank/n910 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[772] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__5_  ( .D(
        \iRF_stage/reg_bank/n911 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[773] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__6_  ( .D(
        \iRF_stage/reg_bank/n912 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[774] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__7_  ( .D(
        \iRF_stage/reg_bank/n913 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[775] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__8_  ( .D(
        \iRF_stage/reg_bank/n914 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[776] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__9_  ( .D(
        \iRF_stage/reg_bank/n915 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[777] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__10_  ( .D(
        \iRF_stage/reg_bank/n916 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[778] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__11_  ( .D(
        \iRF_stage/reg_bank/n917 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[779] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__12_  ( .D(
        \iRF_stage/reg_bank/n918 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[780] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__13_  ( .D(
        \iRF_stage/reg_bank/n919 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[781] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__14_  ( .D(
        \iRF_stage/reg_bank/n920 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[782] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__15_  ( .D(
        \iRF_stage/reg_bank/n921 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[783] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__16_  ( .D(
        \iRF_stage/reg_bank/n922 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[784] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__17_  ( .D(
        \iRF_stage/reg_bank/n923 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[785] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__18_  ( .D(
        \iRF_stage/reg_bank/n924 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[786] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__19_  ( .D(
        \iRF_stage/reg_bank/n925 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[787] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__20_  ( .D(
        \iRF_stage/reg_bank/n926 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[788] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__21_  ( .D(
        \iRF_stage/reg_bank/n927 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[789] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__22_  ( .D(
        \iRF_stage/reg_bank/n928 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[790] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__23_  ( .D(
        \iRF_stage/reg_bank/n929 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[791] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__24_  ( .D(
        \iRF_stage/reg_bank/n930 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[792] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__25_  ( .D(
        \iRF_stage/reg_bank/n931 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[793] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__26_  ( .D(
        \iRF_stage/reg_bank/n932 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[794] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__27_  ( .D(
        \iRF_stage/reg_bank/n933 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[795] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__28_  ( .D(
        \iRF_stage/reg_bank/n934 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[796] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__29_  ( .D(
        \iRF_stage/reg_bank/n935 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[797] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__30_  ( .D(
        \iRF_stage/reg_bank/n936 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[798] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_7__31_  ( .D(
        \iRF_stage/reg_bank/n937 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[799] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__0_  ( .D(
        \iRF_stage/reg_bank/n1034 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[896] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__1_  ( .D(
        \iRF_stage/reg_bank/n1035 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[897] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__2_  ( .D(
        \iRF_stage/reg_bank/n1036 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[898] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__3_  ( .D(
        \iRF_stage/reg_bank/n1037 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[899] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__4_  ( .D(
        \iRF_stage/reg_bank/n1038 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[900] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__5_  ( .D(
        \iRF_stage/reg_bank/n1039 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[901] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__6_  ( .D(
        \iRF_stage/reg_bank/n1040 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[902] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__7_  ( .D(
        \iRF_stage/reg_bank/n1041 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[903] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__8_  ( .D(
        \iRF_stage/reg_bank/n1042 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[904] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__9_  ( .D(
        \iRF_stage/reg_bank/n1043 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[905] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__10_  ( .D(
        \iRF_stage/reg_bank/n1044 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[906] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__11_  ( .D(
        \iRF_stage/reg_bank/n1045 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[907] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__12_  ( .D(
        \iRF_stage/reg_bank/n1046 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[908] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__13_  ( .D(
        \iRF_stage/reg_bank/n1047 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[909] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__14_  ( .D(
        \iRF_stage/reg_bank/n1048 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[910] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__15_  ( .D(
        \iRF_stage/reg_bank/n1049 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[911] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__16_  ( .D(
        \iRF_stage/reg_bank/n1050 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[912] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__17_  ( .D(
        \iRF_stage/reg_bank/n1051 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[913] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__18_  ( .D(
        \iRF_stage/reg_bank/n1052 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[914] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__19_  ( .D(
        \iRF_stage/reg_bank/n1053 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[915] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__20_  ( .D(
        \iRF_stage/reg_bank/n1054 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[916] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__21_  ( .D(
        \iRF_stage/reg_bank/n1055 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[917] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__22_  ( .D(
        \iRF_stage/reg_bank/n1056 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[918] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__23_  ( .D(
        \iRF_stage/reg_bank/n1057 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[919] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__24_  ( .D(
        \iRF_stage/reg_bank/n1058 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[920] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__25_  ( .D(
        \iRF_stage/reg_bank/n1059 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[921] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__26_  ( .D(
        \iRF_stage/reg_bank/n1060 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[922] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__27_  ( .D(
        \iRF_stage/reg_bank/n1061 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[923] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__28_  ( .D(
        \iRF_stage/reg_bank/n1062 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[924] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__29_  ( .D(
        \iRF_stage/reg_bank/n1063 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[925] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__30_  ( .D(
        \iRF_stage/reg_bank/n1064 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[926] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_3__31_  ( .D(
        \iRF_stage/reg_bank/n1065 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[927] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__0_  ( .D(
        \iRF_stage/reg_bank/n170 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[32] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__1_  ( .D(
        \iRF_stage/reg_bank/n171 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[33] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__2_  ( .D(
        \iRF_stage/reg_bank/n172 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[34] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__3_  ( .D(
        \iRF_stage/reg_bank/n173 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[35] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__4_  ( .D(
        \iRF_stage/reg_bank/n174 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[36] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__5_  ( .D(
        \iRF_stage/reg_bank/n175 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[37] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__6_  ( .D(
        \iRF_stage/reg_bank/n176 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[38] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__7_  ( .D(
        \iRF_stage/reg_bank/n177 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[39] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__8_  ( .D(
        \iRF_stage/reg_bank/n178 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[40] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__9_  ( .D(
        \iRF_stage/reg_bank/n179 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[41] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__10_  ( .D(
        \iRF_stage/reg_bank/n180 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[42] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__11_  ( .D(
        \iRF_stage/reg_bank/n181 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[43] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__12_  ( .D(
        \iRF_stage/reg_bank/n182 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[44] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__13_  ( .D(
        \iRF_stage/reg_bank/n183 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[45] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__14_  ( .D(
        \iRF_stage/reg_bank/n184 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[46] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__15_  ( .D(
        \iRF_stage/reg_bank/n185 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[47] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__16_  ( .D(
        \iRF_stage/reg_bank/n186 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[48] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__17_  ( .D(
        \iRF_stage/reg_bank/n187 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[49] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__18_  ( .D(
        \iRF_stage/reg_bank/n188 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[50] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__19_  ( .D(
        \iRF_stage/reg_bank/n189 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[51] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__20_  ( .D(
        \iRF_stage/reg_bank/n190 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[52] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__21_  ( .D(
        \iRF_stage/reg_bank/n191 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[53] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__22_  ( .D(
        \iRF_stage/reg_bank/n192 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[54] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__23_  ( .D(
        \iRF_stage/reg_bank/n193 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[55] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__24_  ( .D(
        \iRF_stage/reg_bank/n194 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[56] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__25_  ( .D(
        \iRF_stage/reg_bank/n195 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[57] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__26_  ( .D(
        \iRF_stage/reg_bank/n196 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[58] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__27_  ( .D(
        \iRF_stage/reg_bank/n197 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[59] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__28_  ( .D(
        \iRF_stage/reg_bank/n198 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[60] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__29_  ( .D(
        \iRF_stage/reg_bank/n199 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[61] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__30_  ( .D(
        \iRF_stage/reg_bank/n200 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[62] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_30__31_  ( .D(
        \iRF_stage/reg_bank/n201 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[63] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__0_  ( .D(
        \iRF_stage/reg_bank/n298 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[160] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__1_  ( .D(
        \iRF_stage/reg_bank/n299 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[161] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__2_  ( .D(
        \iRF_stage/reg_bank/n300 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[162] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__3_  ( .D(
        \iRF_stage/reg_bank/n301 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[163] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__4_  ( .D(
        \iRF_stage/reg_bank/n302 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[164] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__5_  ( .D(
        \iRF_stage/reg_bank/n303 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[165] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__6_  ( .D(
        \iRF_stage/reg_bank/n304 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[166] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__7_  ( .D(
        \iRF_stage/reg_bank/n305 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[167] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__8_  ( .D(
        \iRF_stage/reg_bank/n306 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[168] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__9_  ( .D(
        \iRF_stage/reg_bank/n307 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[169] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__10_  ( .D(
        \iRF_stage/reg_bank/n308 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[170] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__11_  ( .D(
        \iRF_stage/reg_bank/n309 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[171] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__12_  ( .D(
        \iRF_stage/reg_bank/n310 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[172] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__13_  ( .D(
        \iRF_stage/reg_bank/n311 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[173] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__14_  ( .D(
        \iRF_stage/reg_bank/n312 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[174] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__15_  ( .D(
        \iRF_stage/reg_bank/n313 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[175] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__16_  ( .D(
        \iRF_stage/reg_bank/n314 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[176] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__17_  ( .D(
        \iRF_stage/reg_bank/n315 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[177] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__18_  ( .D(
        \iRF_stage/reg_bank/n316 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[178] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__19_  ( .D(
        \iRF_stage/reg_bank/n317 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[179] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__20_  ( .D(
        \iRF_stage/reg_bank/n318 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[180] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__21_  ( .D(
        \iRF_stage/reg_bank/n319 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[181] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__22_  ( .D(
        \iRF_stage/reg_bank/n320 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[182] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__23_  ( .D(
        \iRF_stage/reg_bank/n321 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[183] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__24_  ( .D(
        \iRF_stage/reg_bank/n322 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[184] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__25_  ( .D(
        \iRF_stage/reg_bank/n323 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[185] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__26_  ( .D(
        \iRF_stage/reg_bank/n324 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[186] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__27_  ( .D(
        \iRF_stage/reg_bank/n325 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[187] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__28_  ( .D(
        \iRF_stage/reg_bank/n326 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[188] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__29_  ( .D(
        \iRF_stage/reg_bank/n327 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[189] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__30_  ( .D(
        \iRF_stage/reg_bank/n328 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[190] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_26__31_  ( .D(
        \iRF_stage/reg_bank/n329 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[191] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__0_  ( .D(
        \iRF_stage/reg_bank/n426 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[288] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__1_  ( .D(
        \iRF_stage/reg_bank/n427 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[289] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__2_  ( .D(
        \iRF_stage/reg_bank/n428 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[290] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__3_  ( .D(
        \iRF_stage/reg_bank/n429 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[291] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__4_  ( .D(
        \iRF_stage/reg_bank/n430 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[292] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__5_  ( .D(
        \iRF_stage/reg_bank/n431 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[293] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__6_  ( .D(
        \iRF_stage/reg_bank/n432 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[294] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__7_  ( .D(
        \iRF_stage/reg_bank/n433 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[295] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__8_  ( .D(
        \iRF_stage/reg_bank/n434 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[296] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__9_  ( .D(
        \iRF_stage/reg_bank/n435 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[297] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__10_  ( .D(
        \iRF_stage/reg_bank/n436 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[298] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__11_  ( .D(
        \iRF_stage/reg_bank/n437 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[299] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__12_  ( .D(
        \iRF_stage/reg_bank/n438 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[300] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__13_  ( .D(
        \iRF_stage/reg_bank/n439 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[301] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__14_  ( .D(
        \iRF_stage/reg_bank/n440 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[302] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__15_  ( .D(
        \iRF_stage/reg_bank/n441 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[303] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__16_  ( .D(
        \iRF_stage/reg_bank/n442 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[304] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__17_  ( .D(
        \iRF_stage/reg_bank/n443 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[305] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__18_  ( .D(
        \iRF_stage/reg_bank/n444 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[306] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__19_  ( .D(
        \iRF_stage/reg_bank/n445 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[307] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__20_  ( .D(
        \iRF_stage/reg_bank/n446 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[308] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__21_  ( .D(
        \iRF_stage/reg_bank/n447 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[309] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__22_  ( .D(
        \iRF_stage/reg_bank/n448 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[310] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__23_  ( .D(
        \iRF_stage/reg_bank/n449 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[311] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__24_  ( .D(
        \iRF_stage/reg_bank/n450 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[312] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__25_  ( .D(
        \iRF_stage/reg_bank/n451 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[313] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__26_  ( .D(
        \iRF_stage/reg_bank/n452 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[314] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__27_  ( .D(
        \iRF_stage/reg_bank/n453 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[315] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__28_  ( .D(
        \iRF_stage/reg_bank/n454 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[316] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__29_  ( .D(
        \iRF_stage/reg_bank/n455 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[317] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__30_  ( .D(
        \iRF_stage/reg_bank/n456 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[318] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_22__31_  ( .D(
        \iRF_stage/reg_bank/n457 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[319] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__0_  ( .D(
        \iRF_stage/reg_bank/n554 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[416] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__1_  ( .D(
        \iRF_stage/reg_bank/n555 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[417] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__2_  ( .D(
        \iRF_stage/reg_bank/n556 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[418] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__3_  ( .D(
        \iRF_stage/reg_bank/n557 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[419] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__4_  ( .D(
        \iRF_stage/reg_bank/n558 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[420] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__5_  ( .D(
        \iRF_stage/reg_bank/n559 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[421] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__6_  ( .D(
        \iRF_stage/reg_bank/n560 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[422] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__7_  ( .D(
        \iRF_stage/reg_bank/n561 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[423] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__8_  ( .D(
        \iRF_stage/reg_bank/n562 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[424] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__9_  ( .D(
        \iRF_stage/reg_bank/n563 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[425] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__10_  ( .D(
        \iRF_stage/reg_bank/n564 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[426] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__11_  ( .D(
        \iRF_stage/reg_bank/n565 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[427] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__12_  ( .D(
        \iRF_stage/reg_bank/n566 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[428] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__13_  ( .D(
        \iRF_stage/reg_bank/n567 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[429] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__14_  ( .D(
        \iRF_stage/reg_bank/n568 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[430] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__15_  ( .D(
        \iRF_stage/reg_bank/n569 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[431] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__16_  ( .D(
        \iRF_stage/reg_bank/n570 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[432] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__17_  ( .D(
        \iRF_stage/reg_bank/n571 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[433] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__18_  ( .D(
        \iRF_stage/reg_bank/n572 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[434] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__19_  ( .D(
        \iRF_stage/reg_bank/n573 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[435] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__20_  ( .D(
        \iRF_stage/reg_bank/n574 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[436] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__21_  ( .D(
        \iRF_stage/reg_bank/n575 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[437] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__22_  ( .D(
        \iRF_stage/reg_bank/n576 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[438] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__23_  ( .D(
        \iRF_stage/reg_bank/n577 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[439] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__24_  ( .D(
        \iRF_stage/reg_bank/n578 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[440] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__25_  ( .D(
        \iRF_stage/reg_bank/n579 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[441] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__26_  ( .D(
        \iRF_stage/reg_bank/n580 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[442] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__27_  ( .D(
        \iRF_stage/reg_bank/n581 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[443] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__28_  ( .D(
        \iRF_stage/reg_bank/n582 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[444] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__29_  ( .D(
        \iRF_stage/reg_bank/n583 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[445] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__30_  ( .D(
        \iRF_stage/reg_bank/n584 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[446] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_18__31_  ( .D(
        \iRF_stage/reg_bank/n585 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[447] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__0_  ( .D(
        \iRF_stage/reg_bank/n682 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[544] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__1_  ( .D(
        \iRF_stage/reg_bank/n683 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[545] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__2_  ( .D(
        \iRF_stage/reg_bank/n684 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[546] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__3_  ( .D(
        \iRF_stage/reg_bank/n685 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[547] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__4_  ( .D(
        \iRF_stage/reg_bank/n686 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[548] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__5_  ( .D(
        \iRF_stage/reg_bank/n687 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[549] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__6_  ( .D(
        \iRF_stage/reg_bank/n688 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[550] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__7_  ( .D(
        \iRF_stage/reg_bank/n689 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[551] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__8_  ( .D(
        \iRF_stage/reg_bank/n690 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[552] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__9_  ( .D(
        \iRF_stage/reg_bank/n691 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[553] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__10_  ( .D(
        \iRF_stage/reg_bank/n692 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[554] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__11_  ( .D(
        \iRF_stage/reg_bank/n693 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[555] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__12_  ( .D(
        \iRF_stage/reg_bank/n694 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[556] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__13_  ( .D(
        \iRF_stage/reg_bank/n695 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[557] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__14_  ( .D(
        \iRF_stage/reg_bank/n696 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[558] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__15_  ( .D(
        \iRF_stage/reg_bank/n697 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[559] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__16_  ( .D(
        \iRF_stage/reg_bank/n698 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[560] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__17_  ( .D(
        \iRF_stage/reg_bank/n699 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[561] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__18_  ( .D(
        \iRF_stage/reg_bank/n700 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[562] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__19_  ( .D(
        \iRF_stage/reg_bank/n701 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[563] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__20_  ( .D(
        \iRF_stage/reg_bank/n702 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[564] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__21_  ( .D(
        \iRF_stage/reg_bank/n703 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[565] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__22_  ( .D(
        \iRF_stage/reg_bank/n704 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[566] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__23_  ( .D(
        \iRF_stage/reg_bank/n705 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[567] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__24_  ( .D(
        \iRF_stage/reg_bank/n706 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[568] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__25_  ( .D(
        \iRF_stage/reg_bank/n707 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[569] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__26_  ( .D(
        \iRF_stage/reg_bank/n708 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[570] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__27_  ( .D(
        \iRF_stage/reg_bank/n709 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[571] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__28_  ( .D(
        \iRF_stage/reg_bank/n710 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[572] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__29_  ( .D(
        \iRF_stage/reg_bank/n711 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[573] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__30_  ( .D(
        \iRF_stage/reg_bank/n712 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[574] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_14__31_  ( .D(
        \iRF_stage/reg_bank/n713 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[575] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__0_  ( .D(
        \iRF_stage/reg_bank/n810 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[672] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__1_  ( .D(
        \iRF_stage/reg_bank/n811 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[673] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__2_  ( .D(
        \iRF_stage/reg_bank/n812 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[674] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__3_  ( .D(
        \iRF_stage/reg_bank/n813 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[675] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__4_  ( .D(
        \iRF_stage/reg_bank/n814 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[676] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__5_  ( .D(
        \iRF_stage/reg_bank/n815 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[677] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__6_  ( .D(
        \iRF_stage/reg_bank/n816 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[678] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__7_  ( .D(
        \iRF_stage/reg_bank/n817 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[679] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__8_  ( .D(
        \iRF_stage/reg_bank/n818 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[680] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__9_  ( .D(
        \iRF_stage/reg_bank/n819 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[681] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__10_  ( .D(
        \iRF_stage/reg_bank/n820 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[682] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__11_  ( .D(
        \iRF_stage/reg_bank/n821 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[683] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__12_  ( .D(
        \iRF_stage/reg_bank/n822 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[684] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__13_  ( .D(
        \iRF_stage/reg_bank/n823 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[685] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__14_  ( .D(
        \iRF_stage/reg_bank/n824 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[686] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__15_  ( .D(
        \iRF_stage/reg_bank/n825 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[687] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__16_  ( .D(
        \iRF_stage/reg_bank/n826 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[688] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__17_  ( .D(
        \iRF_stage/reg_bank/n827 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[689] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__18_  ( .D(
        \iRF_stage/reg_bank/n828 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[690] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__19_  ( .D(
        \iRF_stage/reg_bank/n829 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[691] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__20_  ( .D(
        \iRF_stage/reg_bank/n830 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[692] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__21_  ( .D(
        \iRF_stage/reg_bank/n831 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[693] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__22_  ( .D(
        \iRF_stage/reg_bank/n832 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[694] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__23_  ( .D(
        \iRF_stage/reg_bank/n833 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[695] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__24_  ( .D(
        \iRF_stage/reg_bank/n834 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[696] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__25_  ( .D(
        \iRF_stage/reg_bank/n835 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[697] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__26_  ( .D(
        \iRF_stage/reg_bank/n836 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[698] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__27_  ( .D(
        \iRF_stage/reg_bank/n837 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[699] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__28_  ( .D(
        \iRF_stage/reg_bank/n838 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[700] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__29_  ( .D(
        \iRF_stage/reg_bank/n839 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[701] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__30_  ( .D(
        \iRF_stage/reg_bank/n840 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[702] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_10__31_  ( .D(
        \iRF_stage/reg_bank/n841 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[703] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__0_  ( .D(
        \iRF_stage/reg_bank/n938 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[800] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__1_  ( .D(
        \iRF_stage/reg_bank/n939 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[801] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__2_  ( .D(
        \iRF_stage/reg_bank/n940 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[802] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__3_  ( .D(
        \iRF_stage/reg_bank/n941 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[803] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__4_  ( .D(
        \iRF_stage/reg_bank/n942 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[804] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__5_  ( .D(
        \iRF_stage/reg_bank/n943 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[805] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__6_  ( .D(
        \iRF_stage/reg_bank/n944 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[806] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__7_  ( .D(
        \iRF_stage/reg_bank/n945 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[807] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__8_  ( .D(
        \iRF_stage/reg_bank/n946 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[808] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__9_  ( .D(
        \iRF_stage/reg_bank/n947 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[809] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__10_  ( .D(
        \iRF_stage/reg_bank/n948 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[810] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__11_  ( .D(
        \iRF_stage/reg_bank/n949 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[811] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__12_  ( .D(
        \iRF_stage/reg_bank/n950 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[812] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__13_  ( .D(
        \iRF_stage/reg_bank/n951 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[813] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__14_  ( .D(
        \iRF_stage/reg_bank/n952 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[814] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__15_  ( .D(
        \iRF_stage/reg_bank/n953 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[815] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__16_  ( .D(
        \iRF_stage/reg_bank/n954 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[816] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__17_  ( .D(
        \iRF_stage/reg_bank/n955 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[817] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__18_  ( .D(
        \iRF_stage/reg_bank/n956 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[818] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__19_  ( .D(
        \iRF_stage/reg_bank/n957 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[819] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__20_  ( .D(
        \iRF_stage/reg_bank/n958 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[820] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__21_  ( .D(
        \iRF_stage/reg_bank/n959 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[821] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__22_  ( .D(
        \iRF_stage/reg_bank/n960 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[822] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__23_  ( .D(
        \iRF_stage/reg_bank/n961 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[823] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__24_  ( .D(
        \iRF_stage/reg_bank/n962 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[824] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__25_  ( .D(
        \iRF_stage/reg_bank/n963 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[825] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__26_  ( .D(
        \iRF_stage/reg_bank/n964 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[826] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__27_  ( .D(
        \iRF_stage/reg_bank/n965 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[827] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__28_  ( .D(
        \iRF_stage/reg_bank/n966 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[828] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__29_  ( .D(
        \iRF_stage/reg_bank/n967 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[829] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__30_  ( .D(
        \iRF_stage/reg_bank/n968 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[830] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_6__31_  ( .D(
        \iRF_stage/reg_bank/n969 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[831] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__0_  ( .D(
        \iRF_stage/reg_bank/n1066 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[928] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__1_  ( .D(
        \iRF_stage/reg_bank/n1067 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[929] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__2_  ( .D(
        \iRF_stage/reg_bank/n1068 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[930] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__3_  ( .D(
        \iRF_stage/reg_bank/n1069 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[931] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__4_  ( .D(
        \iRF_stage/reg_bank/n1070 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[932] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__5_  ( .D(
        \iRF_stage/reg_bank/n1071 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[933] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__6_  ( .D(
        \iRF_stage/reg_bank/n1072 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[934] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__7_  ( .D(
        \iRF_stage/reg_bank/n1073 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[935] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__8_  ( .D(
        \iRF_stage/reg_bank/n1074 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[936] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__9_  ( .D(
        \iRF_stage/reg_bank/n1075 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[937] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__10_  ( .D(
        \iRF_stage/reg_bank/n1076 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[938] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__11_  ( .D(
        \iRF_stage/reg_bank/n1077 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[939] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__12_  ( .D(
        \iRF_stage/reg_bank/n1078 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[940] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__13_  ( .D(
        \iRF_stage/reg_bank/n1079 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[941] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__14_  ( .D(
        \iRF_stage/reg_bank/n1080 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[942] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__15_  ( .D(
        \iRF_stage/reg_bank/n1081 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[943] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__16_  ( .D(
        \iRF_stage/reg_bank/n1082 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[944] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__17_  ( .D(
        \iRF_stage/reg_bank/n1083 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[945] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__18_  ( .D(
        \iRF_stage/reg_bank/n1084 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[946] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__19_  ( .D(
        \iRF_stage/reg_bank/n1085 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[947] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__20_  ( .D(
        \iRF_stage/reg_bank/n1086 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[948] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__21_  ( .D(
        \iRF_stage/reg_bank/n1087 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[949] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__22_  ( .D(
        \iRF_stage/reg_bank/n1088 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[950] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__23_  ( .D(
        \iRF_stage/reg_bank/n1089 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[951] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__24_  ( .D(
        \iRF_stage/reg_bank/n1090 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[952] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__25_  ( .D(
        \iRF_stage/reg_bank/n1091 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[953] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__26_  ( .D(
        \iRF_stage/reg_bank/n1092 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[954] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__27_  ( .D(
        \iRF_stage/reg_bank/n1093 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[955] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__28_  ( .D(
        \iRF_stage/reg_bank/n1094 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[956] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__29_  ( .D(
        \iRF_stage/reg_bank/n1095 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[957] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__30_  ( .D(
        \iRF_stage/reg_bank/n1096 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[958] ) );
  DFFHQX1 \iRF_stage/reg_bank/reg_bank_reg_2__31_  ( .D(
        \iRF_stage/reg_bank/n1097 ), .CK(clk), .Q(
        \iRF_stage/reg_bank/reg_bank[959] ) );
  DFFHQX1 \rnd_pass2/r5_o_reg_0_  ( .D(BUS1724[0]), .CK(clk), .Q(BUS18211[0])
         );
  DFFHQX1 \iRF_stage/reg_bank/r_wraddress_reg_3_  ( .D(BUS18211[3]), .CK(clk), 
        .Q(\iRF_stage/reg_bank/r_wraddress[3] ) );
  DFFHQX1 \iRF_stage/reg_bank/r_wren_reg  ( .D(NET1375), .CK(clk), .Q(
        \iRF_stage/reg_bank/r_wren ) );
  DFFHQX1 \rnd_pass2/r5_o_reg_1_  ( .D(BUS1724[1]), .CK(clk), .Q(BUS18211[1])
         );
  DFFTRX1 \iRF_stage/MAIN_FSM/delay_counter_reg_0_  ( .D(n1937), .RN(
        \iRF_stage/MAIN_FSM/n57 ), .CK(clk), .Q(
        \iRF_stage/MAIN_FSM/delay_counter[0] ), .QN(n1937) );
  DFFHQX1 \iRF_stage/reg_bank/r_wraddress_reg_0_  ( .D(BUS18211[0]), .CK(clk), 
        .Q(\iRF_stage/reg_bank/r_wraddress[0] ) );
  DFFHQX1 \iRF_stage/MAIN_FSM/CurrState_reg_2_  ( .D(\iRF_stage/MAIN_FSM/N52 ), 
        .CK(clk), .Q(\iRF_stage/MAIN_FSM/CurrState[2] ) );
  DFFHQX1 \pc/r32_o_reg_0_  ( .D(pc_o[0]), .CK(clk), .Q(
        \iRF_stage/i_pc_gen/N34 ) );
  DFFHQX1 \pc/r32_o_reg_1_  ( .D(pc_o[1]), .CK(clk), .Q(BUS27031[1]) );
  DFFHQX1 \rnd_pass1/r5_o_reg_4_  ( .D(BUS1726[4]), .CK(clk), .Q(BUS1724[4])
         );
  DFFHQX1 \iRF_stage/MAIN_FSM/CurrState_reg_0_  ( .D(\iRF_stage/MAIN_FSM/N50 ), 
        .CK(clk), .Q(\iRF_stage/MAIN_FSM/CurrState[0] ) );
  DFFHQX1 \rnd_pass2/r5_o_reg_2_  ( .D(BUS1724[2]), .CK(clk), .Q(BUS18211[2])
         );
  DFFHQX1 \rnd_pass2/r5_o_reg_3_  ( .D(BUS1724[3]), .CK(clk), .Q(BUS18211[3])
         );
  DFFHQX1 \iRF_stage/reg_bank/r_wraddress_reg_1_  ( .D(BUS18211[1]), .CK(clk), 
        .Q(\iRF_stage/reg_bank/r_wraddress[1] ) );
  DFFHQX1 \iRF_stage/MAIN_FSM/CurrState_reg_1_  ( .D(\iRF_stage/MAIN_FSM/N51 ), 
        .CK(clk), .Q(\iRF_stage/MAIN_FSM/CurrState[1] ) );
  DFFHQX1 \MEM_CTL/dmem_ctl_post/byte_addr_o_reg_1_  ( .D(addr_o[1]), .CK(clk), 
        .Q(\MEM_CTL/BUS629[1] ) );
  DFFHQX1 \rnd_pass1/r5_o_reg_2_  ( .D(BUS1726[2]), .CK(clk), .Q(BUS1724[2])
         );
  DFFHQX1 \rnd_pass1/r5_o_reg_3_  ( .D(BUS1726[3]), .CK(clk), .Q(BUS1724[3])
         );
  DFFHQX1 \iRF_stage/reg_bank/r_wraddress_reg_2_  ( .D(BUS18211[2]), .CK(clk), 
        .Q(\iRF_stage/reg_bank/r_wraddress[2] ) );
  DFFTRX1 \iRF_stage/MAIN_FSM/delay_counter_reg_4_  ( .D(
        \iRF_stage/MAIN_FSM/N36 ), .RN(\iRF_stage/MAIN_FSM/n57 ), .CK(clk), 
        .Q(\iRF_stage/MAIN_FSM/delay_counter[4] ), .QN(n306) );
  DFFHQX1 \pc/r32_o_reg_2_  ( .D(pc_o[2]), .CK(clk), .Q(BUS27031[2]) );
  DFFHQX1 \pc/r32_o_reg_3_  ( .D(pc_o[3]), .CK(clk), .Q(BUS27031[3]) );
  DFFHQX1 \pc/r32_o_reg_4_  ( .D(pc_o[4]), .CK(clk), .Q(BUS27031[4]) );
  DFFHQX1 \pc/r32_o_reg_5_  ( .D(pc_o[5]), .CK(clk), .Q(BUS27031[5]) );
  DFFHQX1 \pc/r32_o_reg_6_  ( .D(pc_o[6]), .CK(clk), .Q(BUS27031[6]) );
  DFFHQX1 \pc/r32_o_reg_7_  ( .D(pc_o[7]), .CK(clk), .Q(BUS27031[7]) );
  DFFHQX1 \pc/r32_o_reg_8_  ( .D(pc_o[8]), .CK(clk), .Q(BUS27031[8]) );
  DFFHQX1 \pc/r32_o_reg_9_  ( .D(pc_o[9]), .CK(clk), .Q(BUS27031[9]) );
  DFFHQX1 \pc/r32_o_reg_10_  ( .D(pc_o[10]), .CK(clk), .Q(BUS27031[10]) );
  DFFHQX1 \pc/r32_o_reg_11_  ( .D(pc_o[11]), .CK(clk), .Q(BUS27031[11]) );
  DFFHQX1 \pc/r32_o_reg_12_  ( .D(pc_o[12]), .CK(clk), .Q(BUS27031[12]) );
  DFFHQX1 \pc/r32_o_reg_13_  ( .D(pc_o[13]), .CK(clk), .Q(BUS27031[13]) );
  DFFHQX1 \pc/r32_o_reg_14_  ( .D(pc_o[14]), .CK(clk), .Q(BUS27031[14]) );
  DFFHQX1 \pc/r32_o_reg_15_  ( .D(pc_o[15]), .CK(clk), .Q(BUS27031[15]) );
  DFFHQX1 \pc/r32_o_reg_16_  ( .D(pc_o[16]), .CK(clk), .Q(BUS27031[16]) );
  DFFHQX1 \pc/r32_o_reg_17_  ( .D(pc_o[17]), .CK(clk), .Q(BUS27031[17]) );
  DFFHQX1 \pc/r32_o_reg_18_  ( .D(pc_o[18]), .CK(clk), .Q(BUS27031[18]) );
  DFFHQX1 \pc/r32_o_reg_19_  ( .D(pc_o[19]), .CK(clk), .Q(BUS27031[19]) );
  DFFHQX1 \pc/r32_o_reg_20_  ( .D(pc_o[20]), .CK(clk), .Q(BUS27031[20]) );
  DFFHQX1 \pc/r32_o_reg_21_  ( .D(pc_o[21]), .CK(clk), .Q(BUS27031[21]) );
  DFFHQX1 \pc/r32_o_reg_22_  ( .D(pc_o[22]), .CK(clk), .Q(BUS27031[22]) );
  DFFHQX1 \pc/r32_o_reg_23_  ( .D(pc_o[23]), .CK(clk), .Q(BUS27031[23]) );
  DFFHQX1 \pc/r32_o_reg_24_  ( .D(pc_o[24]), .CK(clk), .Q(BUS27031[24]) );
  DFFHQX1 \pc/r32_o_reg_25_  ( .D(pc_o[25]), .CK(clk), .Q(BUS27031[25]) );
  DFFHQX1 \pc/r32_o_reg_26_  ( .D(pc_o[26]), .CK(clk), .Q(BUS27031[26]) );
  DFFHQX1 \pc/r32_o_reg_27_  ( .D(pc_o[27]), .CK(clk), .Q(BUS27031[27]) );
  DFFHQX1 \pc/r32_o_reg_28_  ( .D(pc_o[28]), .CK(clk), .Q(BUS27031[28]) );
  DFFHQX1 \pc/r32_o_reg_29_  ( .D(pc_o[29]), .CK(clk), .Q(BUS27031[29]) );
  DFFHQX1 \pc/r32_o_reg_30_  ( .D(pc_o[30]), .CK(clk), .Q(BUS27031[30]) );
  DFFHQX1 \pc/r32_o_reg_31_  ( .D(pc_o[31]), .CK(clk), .Q(BUS27031[31]) );
  DFFTRX1 \iRF_stage/MAIN_FSM/delay_counter_reg_2_  ( .D(
        \iRF_stage/MAIN_FSM/N34 ), .RN(\iRF_stage/MAIN_FSM/n57 ), .CK(clk), 
        .Q(\iRF_stage/MAIN_FSM/delay_counter[2] ) );
  DFFTRX1 \iRF_stage/MAIN_FSM/delay_counter_reg_3_  ( .D(
        \iRF_stage/MAIN_FSM/N35 ), .RN(\iRF_stage/MAIN_FSM/n57 ), .CK(clk), 
        .Q(\iRF_stage/MAIN_FSM/delay_counter[3] ) );
  DFFTRX1 \iRF_stage/MAIN_FSM/delay_counter_reg_1_  ( .D(
        \iRF_stage/MAIN_FSM/N33 ), .RN(\iRF_stage/MAIN_FSM/n57 ), .CK(clk), 
        .Q(\iRF_stage/MAIN_FSM/delay_counter[1] ) );
  EDFFX1 \iRF_stage/reg_bank/r_rdaddress_b_reg_0_  ( .D(\iRF_stage/BUS3236[0] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N17 ), .QN(n339) );
  EDFFX1 \iRF_stage/reg_bank/r_rdaddress_b_reg_1_  ( .D(\iRF_stage/BUS3236[1] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N18 ), .QN(n340) );
  EDFFX1 \iRF_stage/reg_bank/r_rdaddress_a_reg_0_  ( .D(\iRF_stage/BUS3237[0] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N12 ), .QN(n334) );
  EDFFX1 \iRF_stage/reg_bank/r_rdaddress_a_reg_1_  ( .D(\iRF_stage/BUS3237[1] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N13 ), .QN(n335) );
  DFFHQX1 \decoder_pipe/pipereg/U18/wb_mux_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5790[0] ), .CK(clk), .Q(NET457) );
  EDFFX2 \iRF_stage/reg_bank/r_rdaddress_b_reg_4_  ( .D(\iRF_stage/BUS3236[4] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N21 ), .QN(n333) );
  EDFFX2 \iRF_stage/reg_bank/r_rdaddress_a_reg_4_  ( .D(\iRF_stage/BUS3237[4] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N16 ), .QN(n338) );
  ADDHXL \iRF_stage/MAIN_FSM/add_58/U1_1_4  ( .A(
        \iRF_stage/MAIN_FSM/delay_counter[4] ), .B(
        \iRF_stage/MAIN_FSM/add_58/carry[4] ), .CO(
        \iRF_stage/MAIN_FSM/add_58/carry[5] ), .S(\iRF_stage/MAIN_FSM/N36 ) );
  XOR3X2 \iexec_stage/add4/add_39/U1_31  ( .A(BUS27031[31]), .B(1'b0), .C(
        \iexec_stage/add4/add_39/carry[31] ), .Y(\iexec_stage/BUS2446[31] ) );
  XOR3X2 \iRF_stage/i_pc_gen/add_70/U1_31  ( .A(BUS27031[31]), .B(BUS7219[31]), 
        .C(\iRF_stage/i_pc_gen/add_70/carry[31] ), .Y(
        \iRF_stage/i_pc_gen/br_addr[31] ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_0  ( .A(\iRF_stage/i_pc_gen/N34 ), .B(
        BUS7219[0]), .CI(1'b0), .CO(\iRF_stage/i_pc_gen/add_70/carry[1] ), .S(
        \iRF_stage/i_pc_gen/br_addr[0] ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_1  ( .A(BUS27031[1]), .B(BUS7219[1]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[1] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[2] ), .S(
        \iRF_stage/i_pc_gen/br_addr[1] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_4  ( .A(BUS27031[4]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[4] ), .CO(
        \iexec_stage/add4/add_39/carry[5] ), .S(\iexec_stage/BUS2446[4] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_5  ( .A(BUS27031[5]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[5] ), .CO(
        \iexec_stage/add4/add_39/carry[6] ), .S(\iexec_stage/BUS2446[5] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_6  ( .A(BUS27031[6]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[6] ), .CO(
        \iexec_stage/add4/add_39/carry[7] ), .S(\iexec_stage/BUS2446[6] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_7  ( .A(BUS27031[7]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[7] ), .CO(
        \iexec_stage/add4/add_39/carry[8] ), .S(\iexec_stage/BUS2446[7] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_8  ( .A(BUS27031[8]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[8] ), .CO(
        \iexec_stage/add4/add_39/carry[9] ), .S(\iexec_stage/BUS2446[8] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_9  ( .A(BUS27031[9]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[9] ), .CO(
        \iexec_stage/add4/add_39/carry[10] ), .S(\iexec_stage/BUS2446[9] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_10  ( .A(BUS27031[10]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[10] ), .CO(
        \iexec_stage/add4/add_39/carry[11] ), .S(\iexec_stage/BUS2446[10] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_11  ( .A(BUS27031[11]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[11] ), .CO(
        \iexec_stage/add4/add_39/carry[12] ), .S(\iexec_stage/BUS2446[11] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_12  ( .A(BUS27031[12]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[12] ), .CO(
        \iexec_stage/add4/add_39/carry[13] ), .S(\iexec_stage/BUS2446[12] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_13  ( .A(BUS27031[13]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[13] ), .CO(
        \iexec_stage/add4/add_39/carry[14] ), .S(\iexec_stage/BUS2446[13] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_14  ( .A(BUS27031[14]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[14] ), .CO(
        \iexec_stage/add4/add_39/carry[15] ), .S(\iexec_stage/BUS2446[14] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_15  ( .A(BUS27031[15]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[15] ), .CO(
        \iexec_stage/add4/add_39/carry[16] ), .S(\iexec_stage/BUS2446[15] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_16  ( .A(BUS27031[16]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[16] ), .CO(
        \iexec_stage/add4/add_39/carry[17] ), .S(\iexec_stage/BUS2446[16] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_17  ( .A(BUS27031[17]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[17] ), .CO(
        \iexec_stage/add4/add_39/carry[18] ), .S(\iexec_stage/BUS2446[17] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_18  ( .A(BUS27031[18]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[18] ), .CO(
        \iexec_stage/add4/add_39/carry[19] ), .S(\iexec_stage/BUS2446[18] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_19  ( .A(BUS27031[19]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[19] ), .CO(
        \iexec_stage/add4/add_39/carry[20] ), .S(\iexec_stage/BUS2446[19] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_20  ( .A(BUS27031[20]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[20] ), .CO(
        \iexec_stage/add4/add_39/carry[21] ), .S(\iexec_stage/BUS2446[20] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_21  ( .A(BUS27031[21]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[21] ), .CO(
        \iexec_stage/add4/add_39/carry[22] ), .S(\iexec_stage/BUS2446[21] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_22  ( .A(BUS27031[22]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[22] ), .CO(
        \iexec_stage/add4/add_39/carry[23] ), .S(\iexec_stage/BUS2446[22] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_23  ( .A(BUS27031[23]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[23] ), .CO(
        \iexec_stage/add4/add_39/carry[24] ), .S(\iexec_stage/BUS2446[23] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_24  ( .A(BUS27031[24]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[24] ), .CO(
        \iexec_stage/add4/add_39/carry[25] ), .S(\iexec_stage/BUS2446[24] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_25  ( .A(BUS27031[25]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[25] ), .CO(
        \iexec_stage/add4/add_39/carry[26] ), .S(\iexec_stage/BUS2446[25] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_26  ( .A(BUS27031[26]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[26] ), .CO(
        \iexec_stage/add4/add_39/carry[27] ), .S(\iexec_stage/BUS2446[26] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_27  ( .A(BUS27031[27]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[27] ), .CO(
        \iexec_stage/add4/add_39/carry[28] ), .S(\iexec_stage/BUS2446[27] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_28  ( .A(BUS27031[28]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[28] ), .CO(
        \iexec_stage/add4/add_39/carry[29] ), .S(\iexec_stage/BUS2446[28] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_29  ( .A(BUS27031[29]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[29] ), .CO(
        \iexec_stage/add4/add_39/carry[30] ), .S(\iexec_stage/BUS2446[29] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_30  ( .A(BUS27031[30]), .B(1'b0), .CI(
        \iexec_stage/add4/add_39/carry[30] ), .CO(
        \iexec_stage/add4/add_39/carry[31] ), .S(\iexec_stage/BUS2446[30] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_30  ( .A(BUS27031[30]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[30] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[31] ), .S(\iRF_stage/i_pc_gen/N64 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_30  ( .A(BUS27031[30]), .B(BUS7219[30]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[30] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[31] ), .S(
        \iRF_stage/i_pc_gen/br_addr[30] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_29  ( .A(BUS27031[29]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[29] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[30] ), .S(\iRF_stage/i_pc_gen/N63 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_29  ( .A(BUS27031[29]), .B(BUS7219[29]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[29] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[30] ), .S(
        \iRF_stage/i_pc_gen/br_addr[29] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_28  ( .A(BUS27031[28]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[28] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[29] ), .S(\iRF_stage/i_pc_gen/N62 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_28  ( .A(BUS27031[28]), .B(BUS7219[28]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[28] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[29] ), .S(
        \iRF_stage/i_pc_gen/br_addr[28] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_27  ( .A(BUS27031[27]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[27] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[28] ), .S(\iRF_stage/i_pc_gen/N61 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_27  ( .A(BUS27031[27]), .B(BUS7219[27]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[27] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[28] ), .S(
        \iRF_stage/i_pc_gen/br_addr[27] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_26  ( .A(BUS27031[26]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[26] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[27] ), .S(\iRF_stage/i_pc_gen/N60 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_26  ( .A(BUS27031[26]), .B(BUS7219[26]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[26] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[27] ), .S(
        \iRF_stage/i_pc_gen/br_addr[26] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_25  ( .A(BUS27031[25]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[25] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[26] ), .S(\iRF_stage/i_pc_gen/N59 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_25  ( .A(BUS27031[25]), .B(BUS7219[25]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[25] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[26] ), .S(
        \iRF_stage/i_pc_gen/br_addr[25] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_24  ( .A(BUS27031[24]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[24] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[25] ), .S(\iRF_stage/i_pc_gen/N58 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_24  ( .A(BUS27031[24]), .B(BUS7219[24]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[24] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[25] ), .S(
        \iRF_stage/i_pc_gen/br_addr[24] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_23  ( .A(BUS27031[23]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[23] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[24] ), .S(\iRF_stage/i_pc_gen/N57 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_23  ( .A(BUS27031[23]), .B(BUS7219[23]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[23] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[24] ), .S(
        \iRF_stage/i_pc_gen/br_addr[23] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_22  ( .A(BUS27031[22]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[22] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[23] ), .S(\iRF_stage/i_pc_gen/N56 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_22  ( .A(BUS27031[22]), .B(BUS7219[22]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[22] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[23] ), .S(
        \iRF_stage/i_pc_gen/br_addr[22] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_21  ( .A(BUS27031[21]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[21] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[22] ), .S(\iRF_stage/i_pc_gen/N55 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_21  ( .A(BUS27031[21]), .B(BUS7219[21]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[21] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[22] ), .S(
        \iRF_stage/i_pc_gen/br_addr[21] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_20  ( .A(BUS27031[20]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[20] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[21] ), .S(\iRF_stage/i_pc_gen/N54 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_20  ( .A(BUS27031[20]), .B(BUS7219[20]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[20] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[21] ), .S(
        \iRF_stage/i_pc_gen/br_addr[20] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_19  ( .A(BUS27031[19]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[19] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[20] ), .S(\iRF_stage/i_pc_gen/N53 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_19  ( .A(BUS27031[19]), .B(BUS7219[19]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[19] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[20] ), .S(
        \iRF_stage/i_pc_gen/br_addr[19] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_18  ( .A(BUS27031[18]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[18] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[19] ), .S(\iRF_stage/i_pc_gen/N52 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_18  ( .A(BUS27031[18]), .B(BUS7219[18]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[18] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[19] ), .S(
        \iRF_stage/i_pc_gen/br_addr[18] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_17  ( .A(BUS27031[17]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[17] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[18] ), .S(\iRF_stage/i_pc_gen/N51 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_17  ( .A(BUS27031[17]), .B(BUS7219[17]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[17] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[18] ), .S(
        \iRF_stage/i_pc_gen/br_addr[17] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_16  ( .A(BUS27031[16]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[16] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[17] ), .S(\iRF_stage/i_pc_gen/N50 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_16  ( .A(BUS27031[16]), .B(BUS7219[16]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[16] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[17] ), .S(
        \iRF_stage/i_pc_gen/br_addr[16] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_15  ( .A(BUS27031[15]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[15] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[16] ), .S(\iRF_stage/i_pc_gen/N49 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_15  ( .A(BUS27031[15]), .B(BUS7219[15]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[15] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[16] ), .S(
        \iRF_stage/i_pc_gen/br_addr[15] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_14  ( .A(BUS27031[14]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[14] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[15] ), .S(\iRF_stage/i_pc_gen/N48 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_14  ( .A(BUS27031[14]), .B(BUS7219[14]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[14] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[15] ), .S(
        \iRF_stage/i_pc_gen/br_addr[14] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_13  ( .A(BUS27031[13]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[13] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[14] ), .S(\iRF_stage/i_pc_gen/N47 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_13  ( .A(BUS27031[13]), .B(BUS7219[13]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[13] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[14] ), .S(
        \iRF_stage/i_pc_gen/br_addr[13] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_12  ( .A(BUS27031[12]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[12] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[13] ), .S(\iRF_stage/i_pc_gen/N46 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_12  ( .A(BUS27031[12]), .B(BUS7219[12]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[12] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[13] ), .S(
        \iRF_stage/i_pc_gen/br_addr[12] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_11  ( .A(BUS27031[11]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[11] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[12] ), .S(\iRF_stage/i_pc_gen/N45 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_11  ( .A(BUS27031[11]), .B(BUS7219[11]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[11] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[12] ), .S(
        \iRF_stage/i_pc_gen/br_addr[11] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_10  ( .A(BUS27031[10]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[10] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[11] ), .S(\iRF_stage/i_pc_gen/N44 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_10  ( .A(BUS27031[10]), .B(BUS7219[10]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[10] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[11] ), .S(
        \iRF_stage/i_pc_gen/br_addr[10] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_9  ( .A(BUS27031[9]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[9] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[10] ), .S(\iRF_stage/i_pc_gen/N43 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_9  ( .A(BUS27031[9]), .B(BUS7219[9]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[9] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[10] ), .S(
        \iRF_stage/i_pc_gen/br_addr[9] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_8  ( .A(BUS27031[8]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[8] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[9] ), .S(\iRF_stage/i_pc_gen/N42 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_8  ( .A(BUS27031[8]), .B(BUS7219[8]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[8] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[9] ), .S(
        \iRF_stage/i_pc_gen/br_addr[8] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_7  ( .A(BUS27031[7]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[7] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[8] ), .S(\iRF_stage/i_pc_gen/N41 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_7  ( .A(BUS27031[7]), .B(BUS7219[7]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[7] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[8] ), .S(
        \iRF_stage/i_pc_gen/br_addr[7] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_6  ( .A(BUS27031[6]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[6] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[7] ), .S(\iRF_stage/i_pc_gen/N40 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_6  ( .A(BUS27031[6]), .B(BUS7219[6]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[6] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[7] ), .S(
        \iRF_stage/i_pc_gen/br_addr[6] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_5  ( .A(BUS27031[5]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[5] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[6] ), .S(\iRF_stage/i_pc_gen/N39 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_5  ( .A(BUS27031[5]), .B(BUS7219[5]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[5] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[6] ), .S(
        \iRF_stage/i_pc_gen/br_addr[5] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_4  ( .A(BUS27031[4]), .B(1'b0), .CI(
        \iRF_stage/i_pc_gen/r62/carry[4] ), .CO(
        \iRF_stage/i_pc_gen/r62/carry[5] ), .S(\iRF_stage/i_pc_gen/N38 ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_4  ( .A(BUS27031[4]), .B(BUS7219[4]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[4] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[5] ), .S(
        \iRF_stage/i_pc_gen/br_addr[4] ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_3  ( .A(BUS27031[3]), .B(BUS7219[3]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[3] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[4] ), .S(
        \iRF_stage/i_pc_gen/br_addr[3] ) );
  ADDFX2 \iRF_stage/i_pc_gen/add_70/U1_2  ( .A(BUS27031[2]), .B(BUS7219[2]), 
        .CI(\iRF_stage/i_pc_gen/add_70/carry[2] ), .CO(
        \iRF_stage/i_pc_gen/add_70/carry[3] ), .S(
        \iRF_stage/i_pc_gen/br_addr[2] ) );
  ADDFX2 \iexec_stage/add4/add_39/U1_3  ( .A(BUS27031[3]), .B(1'b0), .CI(
        BUS27031[2]), .CO(\iexec_stage/add4/add_39/carry[4] ), .S(
        \iexec_stage/BUS2446[3] ) );
  ADDFX2 \iRF_stage/i_pc_gen/r62/U1_3  ( .A(BUS27031[3]), .B(1'b0), .CI(
        BUS27031[2]), .CO(\iRF_stage/i_pc_gen/r62/carry[4] ), .S(
        \iRF_stage/i_pc_gen/N37 ) );
  ADDHXL \iRF_stage/MAIN_FSM/add_58/U1_1_2  ( .A(
        \iRF_stage/MAIN_FSM/delay_counter[2] ), .B(
        \iRF_stage/MAIN_FSM/add_58/carry[2] ), .CO(
        \iRF_stage/MAIN_FSM/add_58/carry[3] ), .S(\iRF_stage/MAIN_FSM/N34 ) );
  ADDHXL \iRF_stage/MAIN_FSM/add_58/U1_1_3  ( .A(
        \iRF_stage/MAIN_FSM/delay_counter[3] ), .B(
        \iRF_stage/MAIN_FSM/add_58/carry[3] ), .CO(
        \iRF_stage/MAIN_FSM/add_58/carry[4] ), .S(\iRF_stage/MAIN_FSM/N35 ) );
  ADDHXL \iRF_stage/MAIN_FSM/add_58/U1_1_1  ( .A(
        \iRF_stage/MAIN_FSM/delay_counter[1] ), .B(
        \iRF_stage/MAIN_FSM/delay_counter[0] ), .CO(
        \iRF_stage/MAIN_FSM/add_58/carry[2] ), .S(\iRF_stage/MAIN_FSM/N33 ) );
  MX4X1 \iRF_stage/reg_bank/U1504  ( .A(\iRF_stage/reg_bank/reg_bank[224] ), 
        .B(\iRF_stage/reg_bank/reg_bank[192] ), .C(
        \iRF_stage/reg_bank/reg_bank[160] ), .D(
        \iRF_stage/reg_bank/reg_bank[128] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1483 ) );
  MX4X1 \iRF_stage/reg_bank/U1515  ( .A(\iRF_stage/reg_bank/reg_bank[225] ), 
        .B(\iRF_stage/reg_bank/reg_bank[193] ), .C(
        \iRF_stage/reg_bank/reg_bank[161] ), .D(
        \iRF_stage/reg_bank/reg_bank[129] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1493 ) );
  MX4X1 \iRF_stage/reg_bank/U1526  ( .A(\iRF_stage/reg_bank/reg_bank[226] ), 
        .B(\iRF_stage/reg_bank/reg_bank[194] ), .C(
        \iRF_stage/reg_bank/reg_bank[162] ), .D(
        \iRF_stage/reg_bank/reg_bank[130] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1503 ) );
  MX4X1 \iRF_stage/reg_bank/U1537  ( .A(\iRF_stage/reg_bank/reg_bank[227] ), 
        .B(\iRF_stage/reg_bank/reg_bank[195] ), .C(
        \iRF_stage/reg_bank/reg_bank[163] ), .D(
        \iRF_stage/reg_bank/reg_bank[131] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1513 ) );
  MX4X1 \iRF_stage/reg_bank/U1548  ( .A(\iRF_stage/reg_bank/reg_bank[228] ), 
        .B(\iRF_stage/reg_bank/reg_bank[196] ), .C(
        \iRF_stage/reg_bank/reg_bank[164] ), .D(
        \iRF_stage/reg_bank/reg_bank[132] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1523 ) );
  MX4X1 \iRF_stage/reg_bank/U1559  ( .A(\iRF_stage/reg_bank/reg_bank[229] ), 
        .B(\iRF_stage/reg_bank/reg_bank[197] ), .C(
        \iRF_stage/reg_bank/reg_bank[165] ), .D(
        \iRF_stage/reg_bank/reg_bank[133] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1533 ) );
  MX4X1 \iRF_stage/reg_bank/U1570  ( .A(\iRF_stage/reg_bank/reg_bank[230] ), 
        .B(\iRF_stage/reg_bank/reg_bank[198] ), .C(
        \iRF_stage/reg_bank/reg_bank[166] ), .D(
        \iRF_stage/reg_bank/reg_bank[134] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1543 ) );
  MX4X1 \iRF_stage/reg_bank/U1581  ( .A(\iRF_stage/reg_bank/reg_bank[231] ), 
        .B(\iRF_stage/reg_bank/reg_bank[199] ), .C(
        \iRF_stage/reg_bank/reg_bank[167] ), .D(
        \iRF_stage/reg_bank/reg_bank[135] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1553 ) );
  MX4X1 \iRF_stage/reg_bank/U1592  ( .A(\iRF_stage/reg_bank/reg_bank[232] ), 
        .B(\iRF_stage/reg_bank/reg_bank[200] ), .C(
        \iRF_stage/reg_bank/reg_bank[168] ), .D(
        \iRF_stage/reg_bank/reg_bank[136] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1563 ) );
  MX4X1 \iRF_stage/reg_bank/U1603  ( .A(\iRF_stage/reg_bank/reg_bank[233] ), 
        .B(\iRF_stage/reg_bank/reg_bank[201] ), .C(
        \iRF_stage/reg_bank/reg_bank[169] ), .D(
        \iRF_stage/reg_bank/reg_bank[137] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1573 ) );
  MX4X1 \iRF_stage/reg_bank/U1614  ( .A(\iRF_stage/reg_bank/reg_bank[234] ), 
        .B(\iRF_stage/reg_bank/reg_bank[202] ), .C(
        \iRF_stage/reg_bank/reg_bank[170] ), .D(
        \iRF_stage/reg_bank/reg_bank[138] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1583 ) );
  MX4X1 \iRF_stage/reg_bank/U1625  ( .A(\iRF_stage/reg_bank/reg_bank[235] ), 
        .B(\iRF_stage/reg_bank/reg_bank[203] ), .C(
        \iRF_stage/reg_bank/reg_bank[171] ), .D(
        \iRF_stage/reg_bank/reg_bank[139] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1593 ) );
  MX4X1 \iRF_stage/reg_bank/U1636  ( .A(\iRF_stage/reg_bank/reg_bank[236] ), 
        .B(\iRF_stage/reg_bank/reg_bank[204] ), .C(
        \iRF_stage/reg_bank/reg_bank[172] ), .D(
        \iRF_stage/reg_bank/reg_bank[140] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1603 ) );
  MX4X1 \iRF_stage/reg_bank/U1647  ( .A(\iRF_stage/reg_bank/reg_bank[237] ), 
        .B(\iRF_stage/reg_bank/reg_bank[205] ), .C(
        \iRF_stage/reg_bank/reg_bank[173] ), .D(
        \iRF_stage/reg_bank/reg_bank[141] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1613 ) );
  MX4X1 \iRF_stage/reg_bank/U1658  ( .A(\iRF_stage/reg_bank/reg_bank[238] ), 
        .B(\iRF_stage/reg_bank/reg_bank[206] ), .C(
        \iRF_stage/reg_bank/reg_bank[174] ), .D(
        \iRF_stage/reg_bank/reg_bank[142] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1623 ) );
  MX4X1 \iRF_stage/reg_bank/U1669  ( .A(\iRF_stage/reg_bank/reg_bank[239] ), 
        .B(\iRF_stage/reg_bank/reg_bank[207] ), .C(
        \iRF_stage/reg_bank/reg_bank[175] ), .D(
        \iRF_stage/reg_bank/reg_bank[143] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1633 ) );
  MX4X1 \iRF_stage/reg_bank/U1680  ( .A(\iRF_stage/reg_bank/reg_bank[240] ), 
        .B(\iRF_stage/reg_bank/reg_bank[208] ), .C(
        \iRF_stage/reg_bank/reg_bank[176] ), .D(
        \iRF_stage/reg_bank/reg_bank[144] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1643 ) );
  MX4X1 \iRF_stage/reg_bank/U1691  ( .A(\iRF_stage/reg_bank/reg_bank[241] ), 
        .B(\iRF_stage/reg_bank/reg_bank[209] ), .C(
        \iRF_stage/reg_bank/reg_bank[177] ), .D(
        \iRF_stage/reg_bank/reg_bank[145] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1653 ) );
  MX4X1 \iRF_stage/reg_bank/U1702  ( .A(\iRF_stage/reg_bank/reg_bank[242] ), 
        .B(\iRF_stage/reg_bank/reg_bank[210] ), .C(
        \iRF_stage/reg_bank/reg_bank[178] ), .D(
        \iRF_stage/reg_bank/reg_bank[146] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1663 ) );
  MX4X1 \iRF_stage/reg_bank/U1713  ( .A(\iRF_stage/reg_bank/reg_bank[243] ), 
        .B(\iRF_stage/reg_bank/reg_bank[211] ), .C(
        \iRF_stage/reg_bank/reg_bank[179] ), .D(
        \iRF_stage/reg_bank/reg_bank[147] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1673 ) );
  MX4X1 \iRF_stage/reg_bank/U1724  ( .A(\iRF_stage/reg_bank/reg_bank[244] ), 
        .B(\iRF_stage/reg_bank/reg_bank[212] ), .C(
        \iRF_stage/reg_bank/reg_bank[180] ), .D(
        \iRF_stage/reg_bank/reg_bank[148] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1683 ) );
  MX4X1 \iRF_stage/reg_bank/U1735  ( .A(\iRF_stage/reg_bank/reg_bank[245] ), 
        .B(\iRF_stage/reg_bank/reg_bank[213] ), .C(
        \iRF_stage/reg_bank/reg_bank[181] ), .D(
        \iRF_stage/reg_bank/reg_bank[149] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1693 ) );
  MX4X1 \iRF_stage/reg_bank/U1746  ( .A(\iRF_stage/reg_bank/reg_bank[246] ), 
        .B(\iRF_stage/reg_bank/reg_bank[214] ), .C(
        \iRF_stage/reg_bank/reg_bank[182] ), .D(
        \iRF_stage/reg_bank/reg_bank[150] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1703 ) );
  MX4X1 \iRF_stage/reg_bank/U1757  ( .A(\iRF_stage/reg_bank/reg_bank[247] ), 
        .B(\iRF_stage/reg_bank/reg_bank[215] ), .C(
        \iRF_stage/reg_bank/reg_bank[183] ), .D(
        \iRF_stage/reg_bank/reg_bank[151] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1713 ) );
  MX4X1 \iRF_stage/reg_bank/U1768  ( .A(\iRF_stage/reg_bank/reg_bank[248] ), 
        .B(\iRF_stage/reg_bank/reg_bank[216] ), .C(
        \iRF_stage/reg_bank/reg_bank[184] ), .D(
        \iRF_stage/reg_bank/reg_bank[152] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1723 ) );
  MX4X1 \iRF_stage/reg_bank/U1779  ( .A(\iRF_stage/reg_bank/reg_bank[249] ), 
        .B(\iRF_stage/reg_bank/reg_bank[217] ), .C(
        \iRF_stage/reg_bank/reg_bank[185] ), .D(
        \iRF_stage/reg_bank/reg_bank[153] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1733 ) );
  MX4X1 \iRF_stage/reg_bank/U1790  ( .A(\iRF_stage/reg_bank/reg_bank[250] ), 
        .B(\iRF_stage/reg_bank/reg_bank[218] ), .C(
        \iRF_stage/reg_bank/reg_bank[186] ), .D(
        \iRF_stage/reg_bank/reg_bank[154] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1743 ) );
  MX4X1 \iRF_stage/reg_bank/U1801  ( .A(\iRF_stage/reg_bank/reg_bank[251] ), 
        .B(\iRF_stage/reg_bank/reg_bank[219] ), .C(
        \iRF_stage/reg_bank/reg_bank[187] ), .D(
        \iRF_stage/reg_bank/reg_bank[155] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1753 ) );
  MX4X1 \iRF_stage/reg_bank/U1812  ( .A(\iRF_stage/reg_bank/reg_bank[252] ), 
        .B(\iRF_stage/reg_bank/reg_bank[220] ), .C(
        \iRF_stage/reg_bank/reg_bank[188] ), .D(
        \iRF_stage/reg_bank/reg_bank[156] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1763 ) );
  MX4X1 \iRF_stage/reg_bank/U1823  ( .A(\iRF_stage/reg_bank/reg_bank[253] ), 
        .B(\iRF_stage/reg_bank/reg_bank[221] ), .C(
        \iRF_stage/reg_bank/reg_bank[189] ), .D(
        \iRF_stage/reg_bank/reg_bank[157] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1773 ) );
  MX4X1 \iRF_stage/reg_bank/U1834  ( .A(\iRF_stage/reg_bank/reg_bank[254] ), 
        .B(\iRF_stage/reg_bank/reg_bank[222] ), .C(
        \iRF_stage/reg_bank/reg_bank[190] ), .D(
        \iRF_stage/reg_bank/reg_bank[158] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1783 ) );
  MX4X1 \iRF_stage/reg_bank/U1845  ( .A(\iRF_stage/reg_bank/reg_bank[255] ), 
        .B(\iRF_stage/reg_bank/reg_bank[223] ), .C(
        \iRF_stage/reg_bank/reg_bank[191] ), .D(
        \iRF_stage/reg_bank/reg_bank[159] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1793 ) );
  MX4X1 \iRF_stage/reg_bank/U1152  ( .A(\iRF_stage/reg_bank/reg_bank[224] ), 
        .B(\iRF_stage/reg_bank/reg_bank[192] ), .C(
        \iRF_stage/reg_bank/reg_bank[160] ), .D(
        \iRF_stage/reg_bank/reg_bank[128] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1163 ) );
  MX4X1 \iRF_stage/reg_bank/U1163  ( .A(\iRF_stage/reg_bank/reg_bank[225] ), 
        .B(\iRF_stage/reg_bank/reg_bank[193] ), .C(
        \iRF_stage/reg_bank/reg_bank[161] ), .D(
        \iRF_stage/reg_bank/reg_bank[129] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1173 ) );
  MX4X1 \iRF_stage/reg_bank/U1174  ( .A(\iRF_stage/reg_bank/reg_bank[226] ), 
        .B(\iRF_stage/reg_bank/reg_bank[194] ), .C(
        \iRF_stage/reg_bank/reg_bank[162] ), .D(
        \iRF_stage/reg_bank/reg_bank[130] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1183 ) );
  MX4X1 \iRF_stage/reg_bank/U1185  ( .A(\iRF_stage/reg_bank/reg_bank[227] ), 
        .B(\iRF_stage/reg_bank/reg_bank[195] ), .C(
        \iRF_stage/reg_bank/reg_bank[163] ), .D(
        \iRF_stage/reg_bank/reg_bank[131] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1193 ) );
  MX4X1 \iRF_stage/reg_bank/U1196  ( .A(\iRF_stage/reg_bank/reg_bank[228] ), 
        .B(\iRF_stage/reg_bank/reg_bank[196] ), .C(
        \iRF_stage/reg_bank/reg_bank[164] ), .D(
        \iRF_stage/reg_bank/reg_bank[132] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1203 ) );
  MX4X1 \iRF_stage/reg_bank/U1207  ( .A(\iRF_stage/reg_bank/reg_bank[229] ), 
        .B(\iRF_stage/reg_bank/reg_bank[197] ), .C(
        \iRF_stage/reg_bank/reg_bank[165] ), .D(
        \iRF_stage/reg_bank/reg_bank[133] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1213 ) );
  MX4X1 \iRF_stage/reg_bank/U1218  ( .A(\iRF_stage/reg_bank/reg_bank[230] ), 
        .B(\iRF_stage/reg_bank/reg_bank[198] ), .C(
        \iRF_stage/reg_bank/reg_bank[166] ), .D(
        \iRF_stage/reg_bank/reg_bank[134] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1223 ) );
  MX4X1 \iRF_stage/reg_bank/U1229  ( .A(\iRF_stage/reg_bank/reg_bank[231] ), 
        .B(\iRF_stage/reg_bank/reg_bank[199] ), .C(
        \iRF_stage/reg_bank/reg_bank[167] ), .D(
        \iRF_stage/reg_bank/reg_bank[135] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1233 ) );
  MX4X1 \iRF_stage/reg_bank/U1240  ( .A(\iRF_stage/reg_bank/reg_bank[232] ), 
        .B(\iRF_stage/reg_bank/reg_bank[200] ), .C(
        \iRF_stage/reg_bank/reg_bank[168] ), .D(
        \iRF_stage/reg_bank/reg_bank[136] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1243 ) );
  MX4X1 \iRF_stage/reg_bank/U1251  ( .A(\iRF_stage/reg_bank/reg_bank[233] ), 
        .B(\iRF_stage/reg_bank/reg_bank[201] ), .C(
        \iRF_stage/reg_bank/reg_bank[169] ), .D(
        \iRF_stage/reg_bank/reg_bank[137] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1253 ) );
  MX4X1 \iRF_stage/reg_bank/U1262  ( .A(\iRF_stage/reg_bank/reg_bank[234] ), 
        .B(\iRF_stage/reg_bank/reg_bank[202] ), .C(
        \iRF_stage/reg_bank/reg_bank[170] ), .D(
        \iRF_stage/reg_bank/reg_bank[138] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1263 ) );
  MX4X1 \iRF_stage/reg_bank/U1273  ( .A(\iRF_stage/reg_bank/reg_bank[235] ), 
        .B(\iRF_stage/reg_bank/reg_bank[203] ), .C(
        \iRF_stage/reg_bank/reg_bank[171] ), .D(
        \iRF_stage/reg_bank/reg_bank[139] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1273 ) );
  MX4X1 \iRF_stage/reg_bank/U1284  ( .A(\iRF_stage/reg_bank/reg_bank[236] ), 
        .B(\iRF_stage/reg_bank/reg_bank[204] ), .C(
        \iRF_stage/reg_bank/reg_bank[172] ), .D(
        \iRF_stage/reg_bank/reg_bank[140] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1283 ) );
  MX4X1 \iRF_stage/reg_bank/U1295  ( .A(\iRF_stage/reg_bank/reg_bank[237] ), 
        .B(\iRF_stage/reg_bank/reg_bank[205] ), .C(
        \iRF_stage/reg_bank/reg_bank[173] ), .D(
        \iRF_stage/reg_bank/reg_bank[141] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1293 ) );
  MX4X1 \iRF_stage/reg_bank/U1306  ( .A(\iRF_stage/reg_bank/reg_bank[238] ), 
        .B(\iRF_stage/reg_bank/reg_bank[206] ), .C(
        \iRF_stage/reg_bank/reg_bank[174] ), .D(
        \iRF_stage/reg_bank/reg_bank[142] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1303 ) );
  MX4X1 \iRF_stage/reg_bank/U1317  ( .A(\iRF_stage/reg_bank/reg_bank[239] ), 
        .B(\iRF_stage/reg_bank/reg_bank[207] ), .C(
        \iRF_stage/reg_bank/reg_bank[175] ), .D(
        \iRF_stage/reg_bank/reg_bank[143] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1313 ) );
  MX4X1 \iRF_stage/reg_bank/U1328  ( .A(\iRF_stage/reg_bank/reg_bank[240] ), 
        .B(\iRF_stage/reg_bank/reg_bank[208] ), .C(
        \iRF_stage/reg_bank/reg_bank[176] ), .D(
        \iRF_stage/reg_bank/reg_bank[144] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1323 ) );
  MX4X1 \iRF_stage/reg_bank/U1339  ( .A(\iRF_stage/reg_bank/reg_bank[241] ), 
        .B(\iRF_stage/reg_bank/reg_bank[209] ), .C(
        \iRF_stage/reg_bank/reg_bank[177] ), .D(
        \iRF_stage/reg_bank/reg_bank[145] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1333 ) );
  MX4X1 \iRF_stage/reg_bank/U1350  ( .A(\iRF_stage/reg_bank/reg_bank[242] ), 
        .B(\iRF_stage/reg_bank/reg_bank[210] ), .C(
        \iRF_stage/reg_bank/reg_bank[178] ), .D(
        \iRF_stage/reg_bank/reg_bank[146] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1343 ) );
  MX4X1 \iRF_stage/reg_bank/U1361  ( .A(\iRF_stage/reg_bank/reg_bank[243] ), 
        .B(\iRF_stage/reg_bank/reg_bank[211] ), .C(
        \iRF_stage/reg_bank/reg_bank[179] ), .D(
        \iRF_stage/reg_bank/reg_bank[147] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1353 ) );
  MX4X1 \iRF_stage/reg_bank/U1372  ( .A(\iRF_stage/reg_bank/reg_bank[244] ), 
        .B(\iRF_stage/reg_bank/reg_bank[212] ), .C(
        \iRF_stage/reg_bank/reg_bank[180] ), .D(
        \iRF_stage/reg_bank/reg_bank[148] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1363 ) );
  MX4X1 \iRF_stage/reg_bank/U1383  ( .A(\iRF_stage/reg_bank/reg_bank[245] ), 
        .B(\iRF_stage/reg_bank/reg_bank[213] ), .C(
        \iRF_stage/reg_bank/reg_bank[181] ), .D(
        \iRF_stage/reg_bank/reg_bank[149] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1373 ) );
  MX4X1 \iRF_stage/reg_bank/U1394  ( .A(\iRF_stage/reg_bank/reg_bank[246] ), 
        .B(\iRF_stage/reg_bank/reg_bank[214] ), .C(
        \iRF_stage/reg_bank/reg_bank[182] ), .D(
        \iRF_stage/reg_bank/reg_bank[150] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1383 ) );
  MX4X1 \iRF_stage/reg_bank/U1405  ( .A(\iRF_stage/reg_bank/reg_bank[247] ), 
        .B(\iRF_stage/reg_bank/reg_bank[215] ), .C(
        \iRF_stage/reg_bank/reg_bank[183] ), .D(
        \iRF_stage/reg_bank/reg_bank[151] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1393 ) );
  MX4X1 \iRF_stage/reg_bank/U1416  ( .A(\iRF_stage/reg_bank/reg_bank[248] ), 
        .B(\iRF_stage/reg_bank/reg_bank[216] ), .C(
        \iRF_stage/reg_bank/reg_bank[184] ), .D(
        \iRF_stage/reg_bank/reg_bank[152] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1403 ) );
  MX4X1 \iRF_stage/reg_bank/U1427  ( .A(\iRF_stage/reg_bank/reg_bank[249] ), 
        .B(\iRF_stage/reg_bank/reg_bank[217] ), .C(
        \iRF_stage/reg_bank/reg_bank[185] ), .D(
        \iRF_stage/reg_bank/reg_bank[153] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1413 ) );
  MX4X1 \iRF_stage/reg_bank/U1438  ( .A(\iRF_stage/reg_bank/reg_bank[250] ), 
        .B(\iRF_stage/reg_bank/reg_bank[218] ), .C(
        \iRF_stage/reg_bank/reg_bank[186] ), .D(
        \iRF_stage/reg_bank/reg_bank[154] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1423 ) );
  MX4X1 \iRF_stage/reg_bank/U1449  ( .A(\iRF_stage/reg_bank/reg_bank[251] ), 
        .B(\iRF_stage/reg_bank/reg_bank[219] ), .C(
        \iRF_stage/reg_bank/reg_bank[187] ), .D(
        \iRF_stage/reg_bank/reg_bank[155] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1433 ) );
  MX4X1 \iRF_stage/reg_bank/U1460  ( .A(\iRF_stage/reg_bank/reg_bank[252] ), 
        .B(\iRF_stage/reg_bank/reg_bank[220] ), .C(
        \iRF_stage/reg_bank/reg_bank[188] ), .D(
        \iRF_stage/reg_bank/reg_bank[156] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1443 ) );
  MX4X1 \iRF_stage/reg_bank/U1471  ( .A(\iRF_stage/reg_bank/reg_bank[253] ), 
        .B(\iRF_stage/reg_bank/reg_bank[221] ), .C(
        \iRF_stage/reg_bank/reg_bank[189] ), .D(
        \iRF_stage/reg_bank/reg_bank[157] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1453 ) );
  MX4X1 \iRF_stage/reg_bank/U1482  ( .A(\iRF_stage/reg_bank/reg_bank[254] ), 
        .B(\iRF_stage/reg_bank/reg_bank[222] ), .C(
        \iRF_stage/reg_bank/reg_bank[190] ), .D(
        \iRF_stage/reg_bank/reg_bank[158] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1463 ) );
  MX4X1 \iRF_stage/reg_bank/U1493  ( .A(\iRF_stage/reg_bank/reg_bank[255] ), 
        .B(\iRF_stage/reg_bank/reg_bank[223] ), .C(
        \iRF_stage/reg_bank/reg_bank[191] ), .D(
        \iRF_stage/reg_bank/reg_bank[159] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1473 ) );
  MX4X1 \iRF_stage/reg_bank/U1506  ( .A(\iRF_stage/reg_bank/reg_bank[480] ), 
        .B(\iRF_stage/reg_bank/reg_bank[448] ), .C(
        \iRF_stage/reg_bank/reg_bank[416] ), .D(
        \iRF_stage/reg_bank/reg_bank[384] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1485 ) );
  MX4X1 \iRF_stage/reg_bank/U1517  ( .A(\iRF_stage/reg_bank/reg_bank[481] ), 
        .B(\iRF_stage/reg_bank/reg_bank[449] ), .C(
        \iRF_stage/reg_bank/reg_bank[417] ), .D(
        \iRF_stage/reg_bank/reg_bank[385] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1495 ) );
  MX4X1 \iRF_stage/reg_bank/U1528  ( .A(\iRF_stage/reg_bank/reg_bank[482] ), 
        .B(\iRF_stage/reg_bank/reg_bank[450] ), .C(
        \iRF_stage/reg_bank/reg_bank[418] ), .D(
        \iRF_stage/reg_bank/reg_bank[386] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1505 ) );
  MX4X1 \iRF_stage/reg_bank/U1539  ( .A(\iRF_stage/reg_bank/reg_bank[483] ), 
        .B(\iRF_stage/reg_bank/reg_bank[451] ), .C(
        \iRF_stage/reg_bank/reg_bank[419] ), .D(
        \iRF_stage/reg_bank/reg_bank[387] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1515 ) );
  MX4X1 \iRF_stage/reg_bank/U1550  ( .A(\iRF_stage/reg_bank/reg_bank[484] ), 
        .B(\iRF_stage/reg_bank/reg_bank[452] ), .C(
        \iRF_stage/reg_bank/reg_bank[420] ), .D(
        \iRF_stage/reg_bank/reg_bank[388] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1525 ) );
  MX4X1 \iRF_stage/reg_bank/U1561  ( .A(\iRF_stage/reg_bank/reg_bank[485] ), 
        .B(\iRF_stage/reg_bank/reg_bank[453] ), .C(
        \iRF_stage/reg_bank/reg_bank[421] ), .D(
        \iRF_stage/reg_bank/reg_bank[389] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1535 ) );
  MX4X1 \iRF_stage/reg_bank/U1572  ( .A(\iRF_stage/reg_bank/reg_bank[486] ), 
        .B(\iRF_stage/reg_bank/reg_bank[454] ), .C(
        \iRF_stage/reg_bank/reg_bank[422] ), .D(
        \iRF_stage/reg_bank/reg_bank[390] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1545 ) );
  MX4X1 \iRF_stage/reg_bank/U1583  ( .A(\iRF_stage/reg_bank/reg_bank[487] ), 
        .B(\iRF_stage/reg_bank/reg_bank[455] ), .C(
        \iRF_stage/reg_bank/reg_bank[423] ), .D(
        \iRF_stage/reg_bank/reg_bank[391] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1555 ) );
  MX4X1 \iRF_stage/reg_bank/U1594  ( .A(\iRF_stage/reg_bank/reg_bank[488] ), 
        .B(\iRF_stage/reg_bank/reg_bank[456] ), .C(
        \iRF_stage/reg_bank/reg_bank[424] ), .D(
        \iRF_stage/reg_bank/reg_bank[392] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1565 ) );
  MX4X1 \iRF_stage/reg_bank/U1605  ( .A(\iRF_stage/reg_bank/reg_bank[489] ), 
        .B(\iRF_stage/reg_bank/reg_bank[457] ), .C(
        \iRF_stage/reg_bank/reg_bank[425] ), .D(
        \iRF_stage/reg_bank/reg_bank[393] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1575 ) );
  MX4X1 \iRF_stage/reg_bank/U1616  ( .A(\iRF_stage/reg_bank/reg_bank[490] ), 
        .B(\iRF_stage/reg_bank/reg_bank[458] ), .C(
        \iRF_stage/reg_bank/reg_bank[426] ), .D(
        \iRF_stage/reg_bank/reg_bank[394] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1585 ) );
  MX4X1 \iRF_stage/reg_bank/U1627  ( .A(\iRF_stage/reg_bank/reg_bank[491] ), 
        .B(\iRF_stage/reg_bank/reg_bank[459] ), .C(
        \iRF_stage/reg_bank/reg_bank[427] ), .D(
        \iRF_stage/reg_bank/reg_bank[395] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1595 ) );
  MX4X1 \iRF_stage/reg_bank/U1638  ( .A(\iRF_stage/reg_bank/reg_bank[492] ), 
        .B(\iRF_stage/reg_bank/reg_bank[460] ), .C(
        \iRF_stage/reg_bank/reg_bank[428] ), .D(
        \iRF_stage/reg_bank/reg_bank[396] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1605 ) );
  MX4X1 \iRF_stage/reg_bank/U1649  ( .A(\iRF_stage/reg_bank/reg_bank[493] ), 
        .B(\iRF_stage/reg_bank/reg_bank[461] ), .C(
        \iRF_stage/reg_bank/reg_bank[429] ), .D(
        \iRF_stage/reg_bank/reg_bank[397] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1615 ) );
  MX4X1 \iRF_stage/reg_bank/U1660  ( .A(\iRF_stage/reg_bank/reg_bank[494] ), 
        .B(\iRF_stage/reg_bank/reg_bank[462] ), .C(
        \iRF_stage/reg_bank/reg_bank[430] ), .D(
        \iRF_stage/reg_bank/reg_bank[398] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1625 ) );
  MX4X1 \iRF_stage/reg_bank/U1671  ( .A(\iRF_stage/reg_bank/reg_bank[495] ), 
        .B(\iRF_stage/reg_bank/reg_bank[463] ), .C(
        \iRF_stage/reg_bank/reg_bank[431] ), .D(
        \iRF_stage/reg_bank/reg_bank[399] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1635 ) );
  MX4X1 \iRF_stage/reg_bank/U1682  ( .A(\iRF_stage/reg_bank/reg_bank[496] ), 
        .B(\iRF_stage/reg_bank/reg_bank[464] ), .C(
        \iRF_stage/reg_bank/reg_bank[432] ), .D(
        \iRF_stage/reg_bank/reg_bank[400] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1645 ) );
  MX4X1 \iRF_stage/reg_bank/U1693  ( .A(\iRF_stage/reg_bank/reg_bank[497] ), 
        .B(\iRF_stage/reg_bank/reg_bank[465] ), .C(
        \iRF_stage/reg_bank/reg_bank[433] ), .D(
        \iRF_stage/reg_bank/reg_bank[401] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1655 ) );
  MX4X1 \iRF_stage/reg_bank/U1704  ( .A(\iRF_stage/reg_bank/reg_bank[498] ), 
        .B(\iRF_stage/reg_bank/reg_bank[466] ), .C(
        \iRF_stage/reg_bank/reg_bank[434] ), .D(
        \iRF_stage/reg_bank/reg_bank[402] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1665 ) );
  MX4X1 \iRF_stage/reg_bank/U1715  ( .A(\iRF_stage/reg_bank/reg_bank[499] ), 
        .B(\iRF_stage/reg_bank/reg_bank[467] ), .C(
        \iRF_stage/reg_bank/reg_bank[435] ), .D(
        \iRF_stage/reg_bank/reg_bank[403] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1675 ) );
  MX4X1 \iRF_stage/reg_bank/U1726  ( .A(\iRF_stage/reg_bank/reg_bank[500] ), 
        .B(\iRF_stage/reg_bank/reg_bank[468] ), .C(
        \iRF_stage/reg_bank/reg_bank[436] ), .D(
        \iRF_stage/reg_bank/reg_bank[404] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1685 ) );
  MX4X1 \iRF_stage/reg_bank/U1737  ( .A(\iRF_stage/reg_bank/reg_bank[501] ), 
        .B(\iRF_stage/reg_bank/reg_bank[469] ), .C(
        \iRF_stage/reg_bank/reg_bank[437] ), .D(
        \iRF_stage/reg_bank/reg_bank[405] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1695 ) );
  MX4X1 \iRF_stage/reg_bank/U1748  ( .A(\iRF_stage/reg_bank/reg_bank[502] ), 
        .B(\iRF_stage/reg_bank/reg_bank[470] ), .C(
        \iRF_stage/reg_bank/reg_bank[438] ), .D(
        \iRF_stage/reg_bank/reg_bank[406] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1705 ) );
  MX4X1 \iRF_stage/reg_bank/U1759  ( .A(\iRF_stage/reg_bank/reg_bank[503] ), 
        .B(\iRF_stage/reg_bank/reg_bank[471] ), .C(
        \iRF_stage/reg_bank/reg_bank[439] ), .D(
        \iRF_stage/reg_bank/reg_bank[407] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1715 ) );
  MX4X1 \iRF_stage/reg_bank/U1770  ( .A(\iRF_stage/reg_bank/reg_bank[504] ), 
        .B(\iRF_stage/reg_bank/reg_bank[472] ), .C(
        \iRF_stage/reg_bank/reg_bank[440] ), .D(
        \iRF_stage/reg_bank/reg_bank[408] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1725 ) );
  MX4X1 \iRF_stage/reg_bank/U1781  ( .A(\iRF_stage/reg_bank/reg_bank[505] ), 
        .B(\iRF_stage/reg_bank/reg_bank[473] ), .C(
        \iRF_stage/reg_bank/reg_bank[441] ), .D(
        \iRF_stage/reg_bank/reg_bank[409] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1735 ) );
  MX4X1 \iRF_stage/reg_bank/U1792  ( .A(\iRF_stage/reg_bank/reg_bank[506] ), 
        .B(\iRF_stage/reg_bank/reg_bank[474] ), .C(
        \iRF_stage/reg_bank/reg_bank[442] ), .D(
        \iRF_stage/reg_bank/reg_bank[410] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1745 ) );
  MX4X1 \iRF_stage/reg_bank/U1803  ( .A(\iRF_stage/reg_bank/reg_bank[507] ), 
        .B(\iRF_stage/reg_bank/reg_bank[475] ), .C(
        \iRF_stage/reg_bank/reg_bank[443] ), .D(
        \iRF_stage/reg_bank/reg_bank[411] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1755 ) );
  MX4X1 \iRF_stage/reg_bank/U1814  ( .A(\iRF_stage/reg_bank/reg_bank[508] ), 
        .B(\iRF_stage/reg_bank/reg_bank[476] ), .C(
        \iRF_stage/reg_bank/reg_bank[444] ), .D(
        \iRF_stage/reg_bank/reg_bank[412] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1765 ) );
  MX4X1 \iRF_stage/reg_bank/U1825  ( .A(\iRF_stage/reg_bank/reg_bank[509] ), 
        .B(\iRF_stage/reg_bank/reg_bank[477] ), .C(
        \iRF_stage/reg_bank/reg_bank[445] ), .D(
        \iRF_stage/reg_bank/reg_bank[413] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1775 ) );
  MX4X1 \iRF_stage/reg_bank/U1836  ( .A(\iRF_stage/reg_bank/reg_bank[510] ), 
        .B(\iRF_stage/reg_bank/reg_bank[478] ), .C(
        \iRF_stage/reg_bank/reg_bank[446] ), .D(
        \iRF_stage/reg_bank/reg_bank[414] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1785 ) );
  MX4X1 \iRF_stage/reg_bank/U1847  ( .A(\iRF_stage/reg_bank/reg_bank[511] ), 
        .B(\iRF_stage/reg_bank/reg_bank[479] ), .C(
        \iRF_stage/reg_bank/reg_bank[447] ), .D(
        \iRF_stage/reg_bank/reg_bank[415] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1795 ) );
  MX4X1 \iRF_stage/reg_bank/U1154  ( .A(\iRF_stage/reg_bank/reg_bank[480] ), 
        .B(\iRF_stage/reg_bank/reg_bank[448] ), .C(
        \iRF_stage/reg_bank/reg_bank[416] ), .D(
        \iRF_stage/reg_bank/reg_bank[384] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1165 ) );
  MX4X1 \iRF_stage/reg_bank/U1165  ( .A(\iRF_stage/reg_bank/reg_bank[481] ), 
        .B(\iRF_stage/reg_bank/reg_bank[449] ), .C(
        \iRF_stage/reg_bank/reg_bank[417] ), .D(
        \iRF_stage/reg_bank/reg_bank[385] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1175 ) );
  MX4X1 \iRF_stage/reg_bank/U1176  ( .A(\iRF_stage/reg_bank/reg_bank[482] ), 
        .B(\iRF_stage/reg_bank/reg_bank[450] ), .C(
        \iRF_stage/reg_bank/reg_bank[418] ), .D(
        \iRF_stage/reg_bank/reg_bank[386] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1185 ) );
  MX4X1 \iRF_stage/reg_bank/U1187  ( .A(\iRF_stage/reg_bank/reg_bank[483] ), 
        .B(\iRF_stage/reg_bank/reg_bank[451] ), .C(
        \iRF_stage/reg_bank/reg_bank[419] ), .D(
        \iRF_stage/reg_bank/reg_bank[387] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1195 ) );
  MX4X1 \iRF_stage/reg_bank/U1198  ( .A(\iRF_stage/reg_bank/reg_bank[484] ), 
        .B(\iRF_stage/reg_bank/reg_bank[452] ), .C(
        \iRF_stage/reg_bank/reg_bank[420] ), .D(
        \iRF_stage/reg_bank/reg_bank[388] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1205 ) );
  MX4X1 \iRF_stage/reg_bank/U1209  ( .A(\iRF_stage/reg_bank/reg_bank[485] ), 
        .B(\iRF_stage/reg_bank/reg_bank[453] ), .C(
        \iRF_stage/reg_bank/reg_bank[421] ), .D(
        \iRF_stage/reg_bank/reg_bank[389] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1215 ) );
  MX4X1 \iRF_stage/reg_bank/U1220  ( .A(\iRF_stage/reg_bank/reg_bank[486] ), 
        .B(\iRF_stage/reg_bank/reg_bank[454] ), .C(
        \iRF_stage/reg_bank/reg_bank[422] ), .D(
        \iRF_stage/reg_bank/reg_bank[390] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1225 ) );
  MX4X1 \iRF_stage/reg_bank/U1231  ( .A(\iRF_stage/reg_bank/reg_bank[487] ), 
        .B(\iRF_stage/reg_bank/reg_bank[455] ), .C(
        \iRF_stage/reg_bank/reg_bank[423] ), .D(
        \iRF_stage/reg_bank/reg_bank[391] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1235 ) );
  MX4X1 \iRF_stage/reg_bank/U1242  ( .A(\iRF_stage/reg_bank/reg_bank[488] ), 
        .B(\iRF_stage/reg_bank/reg_bank[456] ), .C(
        \iRF_stage/reg_bank/reg_bank[424] ), .D(
        \iRF_stage/reg_bank/reg_bank[392] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1245 ) );
  MX4X1 \iRF_stage/reg_bank/U1253  ( .A(\iRF_stage/reg_bank/reg_bank[489] ), 
        .B(\iRF_stage/reg_bank/reg_bank[457] ), .C(
        \iRF_stage/reg_bank/reg_bank[425] ), .D(
        \iRF_stage/reg_bank/reg_bank[393] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1255 ) );
  MX4X1 \iRF_stage/reg_bank/U1264  ( .A(\iRF_stage/reg_bank/reg_bank[490] ), 
        .B(\iRF_stage/reg_bank/reg_bank[458] ), .C(
        \iRF_stage/reg_bank/reg_bank[426] ), .D(
        \iRF_stage/reg_bank/reg_bank[394] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1265 ) );
  MX4X1 \iRF_stage/reg_bank/U1275  ( .A(\iRF_stage/reg_bank/reg_bank[491] ), 
        .B(\iRF_stage/reg_bank/reg_bank[459] ), .C(
        \iRF_stage/reg_bank/reg_bank[427] ), .D(
        \iRF_stage/reg_bank/reg_bank[395] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1275 ) );
  MX4X1 \iRF_stage/reg_bank/U1286  ( .A(\iRF_stage/reg_bank/reg_bank[492] ), 
        .B(\iRF_stage/reg_bank/reg_bank[460] ), .C(
        \iRF_stage/reg_bank/reg_bank[428] ), .D(
        \iRF_stage/reg_bank/reg_bank[396] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1285 ) );
  MX4X1 \iRF_stage/reg_bank/U1297  ( .A(\iRF_stage/reg_bank/reg_bank[493] ), 
        .B(\iRF_stage/reg_bank/reg_bank[461] ), .C(
        \iRF_stage/reg_bank/reg_bank[429] ), .D(
        \iRF_stage/reg_bank/reg_bank[397] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1295 ) );
  MX4X1 \iRF_stage/reg_bank/U1308  ( .A(\iRF_stage/reg_bank/reg_bank[494] ), 
        .B(\iRF_stage/reg_bank/reg_bank[462] ), .C(
        \iRF_stage/reg_bank/reg_bank[430] ), .D(
        \iRF_stage/reg_bank/reg_bank[398] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1305 ) );
  MX4X1 \iRF_stage/reg_bank/U1319  ( .A(\iRF_stage/reg_bank/reg_bank[495] ), 
        .B(\iRF_stage/reg_bank/reg_bank[463] ), .C(
        \iRF_stage/reg_bank/reg_bank[431] ), .D(
        \iRF_stage/reg_bank/reg_bank[399] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1315 ) );
  MX4X1 \iRF_stage/reg_bank/U1330  ( .A(\iRF_stage/reg_bank/reg_bank[496] ), 
        .B(\iRF_stage/reg_bank/reg_bank[464] ), .C(
        \iRF_stage/reg_bank/reg_bank[432] ), .D(
        \iRF_stage/reg_bank/reg_bank[400] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1325 ) );
  MX4X1 \iRF_stage/reg_bank/U1341  ( .A(\iRF_stage/reg_bank/reg_bank[497] ), 
        .B(\iRF_stage/reg_bank/reg_bank[465] ), .C(
        \iRF_stage/reg_bank/reg_bank[433] ), .D(
        \iRF_stage/reg_bank/reg_bank[401] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1335 ) );
  MX4X1 \iRF_stage/reg_bank/U1352  ( .A(\iRF_stage/reg_bank/reg_bank[498] ), 
        .B(\iRF_stage/reg_bank/reg_bank[466] ), .C(
        \iRF_stage/reg_bank/reg_bank[434] ), .D(
        \iRF_stage/reg_bank/reg_bank[402] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1345 ) );
  MX4X1 \iRF_stage/reg_bank/U1363  ( .A(\iRF_stage/reg_bank/reg_bank[499] ), 
        .B(\iRF_stage/reg_bank/reg_bank[467] ), .C(
        \iRF_stage/reg_bank/reg_bank[435] ), .D(
        \iRF_stage/reg_bank/reg_bank[403] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1355 ) );
  MX4X1 \iRF_stage/reg_bank/U1374  ( .A(\iRF_stage/reg_bank/reg_bank[500] ), 
        .B(\iRF_stage/reg_bank/reg_bank[468] ), .C(
        \iRF_stage/reg_bank/reg_bank[436] ), .D(
        \iRF_stage/reg_bank/reg_bank[404] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1365 ) );
  MX4X1 \iRF_stage/reg_bank/U1385  ( .A(\iRF_stage/reg_bank/reg_bank[501] ), 
        .B(\iRF_stage/reg_bank/reg_bank[469] ), .C(
        \iRF_stage/reg_bank/reg_bank[437] ), .D(
        \iRF_stage/reg_bank/reg_bank[405] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1375 ) );
  MX4X1 \iRF_stage/reg_bank/U1396  ( .A(\iRF_stage/reg_bank/reg_bank[502] ), 
        .B(\iRF_stage/reg_bank/reg_bank[470] ), .C(
        \iRF_stage/reg_bank/reg_bank[438] ), .D(
        \iRF_stage/reg_bank/reg_bank[406] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1385 ) );
  MX4X1 \iRF_stage/reg_bank/U1407  ( .A(\iRF_stage/reg_bank/reg_bank[503] ), 
        .B(\iRF_stage/reg_bank/reg_bank[471] ), .C(
        \iRF_stage/reg_bank/reg_bank[439] ), .D(
        \iRF_stage/reg_bank/reg_bank[407] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1395 ) );
  MX4X1 \iRF_stage/reg_bank/U1418  ( .A(\iRF_stage/reg_bank/reg_bank[504] ), 
        .B(\iRF_stage/reg_bank/reg_bank[472] ), .C(
        \iRF_stage/reg_bank/reg_bank[440] ), .D(
        \iRF_stage/reg_bank/reg_bank[408] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1405 ) );
  MX4X1 \iRF_stage/reg_bank/U1429  ( .A(\iRF_stage/reg_bank/reg_bank[505] ), 
        .B(\iRF_stage/reg_bank/reg_bank[473] ), .C(
        \iRF_stage/reg_bank/reg_bank[441] ), .D(
        \iRF_stage/reg_bank/reg_bank[409] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1415 ) );
  MX4X1 \iRF_stage/reg_bank/U1440  ( .A(\iRF_stage/reg_bank/reg_bank[506] ), 
        .B(\iRF_stage/reg_bank/reg_bank[474] ), .C(
        \iRF_stage/reg_bank/reg_bank[442] ), .D(
        \iRF_stage/reg_bank/reg_bank[410] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1425 ) );
  MX4X1 \iRF_stage/reg_bank/U1451  ( .A(\iRF_stage/reg_bank/reg_bank[507] ), 
        .B(\iRF_stage/reg_bank/reg_bank[475] ), .C(
        \iRF_stage/reg_bank/reg_bank[443] ), .D(
        \iRF_stage/reg_bank/reg_bank[411] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1435 ) );
  MX4X1 \iRF_stage/reg_bank/U1462  ( .A(\iRF_stage/reg_bank/reg_bank[508] ), 
        .B(\iRF_stage/reg_bank/reg_bank[476] ), .C(
        \iRF_stage/reg_bank/reg_bank[444] ), .D(
        \iRF_stage/reg_bank/reg_bank[412] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1445 ) );
  MX4X1 \iRF_stage/reg_bank/U1473  ( .A(\iRF_stage/reg_bank/reg_bank[509] ), 
        .B(\iRF_stage/reg_bank/reg_bank[477] ), .C(
        \iRF_stage/reg_bank/reg_bank[445] ), .D(
        \iRF_stage/reg_bank/reg_bank[413] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1455 ) );
  MX4X1 \iRF_stage/reg_bank/U1484  ( .A(\iRF_stage/reg_bank/reg_bank[510] ), 
        .B(\iRF_stage/reg_bank/reg_bank[478] ), .C(
        \iRF_stage/reg_bank/reg_bank[446] ), .D(
        \iRF_stage/reg_bank/reg_bank[414] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1465 ) );
  MX4X1 \iRF_stage/reg_bank/U1495  ( .A(\iRF_stage/reg_bank/reg_bank[511] ), 
        .B(\iRF_stage/reg_bank/reg_bank[479] ), .C(
        \iRF_stage/reg_bank/reg_bank[447] ), .D(
        \iRF_stage/reg_bank/reg_bank[415] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1475 ) );
  MX4X1 \iRF_stage/reg_bank/U1503  ( .A(\iRF_stage/reg_bank/reg_bank[96] ), 
        .B(\iRF_stage/reg_bank/reg_bank[64] ), .C(
        \iRF_stage/reg_bank/reg_bank[32] ), .D(
        \iRF_stage/reg_bank/reg_bank[0] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1482 ) );
  MX4X1 \iRF_stage/reg_bank/U1514  ( .A(\iRF_stage/reg_bank/reg_bank[97] ), 
        .B(\iRF_stage/reg_bank/reg_bank[65] ), .C(
        \iRF_stage/reg_bank/reg_bank[33] ), .D(
        \iRF_stage/reg_bank/reg_bank[1] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1492 ) );
  MX4X1 \iRF_stage/reg_bank/U1525  ( .A(\iRF_stage/reg_bank/reg_bank[98] ), 
        .B(\iRF_stage/reg_bank/reg_bank[66] ), .C(
        \iRF_stage/reg_bank/reg_bank[34] ), .D(
        \iRF_stage/reg_bank/reg_bank[2] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1502 ) );
  MX4X1 \iRF_stage/reg_bank/U1536  ( .A(\iRF_stage/reg_bank/reg_bank[99] ), 
        .B(\iRF_stage/reg_bank/reg_bank[67] ), .C(
        \iRF_stage/reg_bank/reg_bank[35] ), .D(
        \iRF_stage/reg_bank/reg_bank[3] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1512 ) );
  MX4X1 \iRF_stage/reg_bank/U1547  ( .A(\iRF_stage/reg_bank/reg_bank[100] ), 
        .B(\iRF_stage/reg_bank/reg_bank[68] ), .C(
        \iRF_stage/reg_bank/reg_bank[36] ), .D(
        \iRF_stage/reg_bank/reg_bank[4] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1522 ) );
  MX4X1 \iRF_stage/reg_bank/U1558  ( .A(\iRF_stage/reg_bank/reg_bank[101] ), 
        .B(\iRF_stage/reg_bank/reg_bank[69] ), .C(
        \iRF_stage/reg_bank/reg_bank[37] ), .D(
        \iRF_stage/reg_bank/reg_bank[5] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1532 ) );
  MX4X1 \iRF_stage/reg_bank/U1569  ( .A(\iRF_stage/reg_bank/reg_bank[102] ), 
        .B(\iRF_stage/reg_bank/reg_bank[70] ), .C(
        \iRF_stage/reg_bank/reg_bank[38] ), .D(
        \iRF_stage/reg_bank/reg_bank[6] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1542 ) );
  MX4X1 \iRF_stage/reg_bank/U1580  ( .A(\iRF_stage/reg_bank/reg_bank[103] ), 
        .B(\iRF_stage/reg_bank/reg_bank[71] ), .C(
        \iRF_stage/reg_bank/reg_bank[39] ), .D(
        \iRF_stage/reg_bank/reg_bank[7] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1552 ) );
  MX4X1 \iRF_stage/reg_bank/U1591  ( .A(\iRF_stage/reg_bank/reg_bank[104] ), 
        .B(\iRF_stage/reg_bank/reg_bank[72] ), .C(
        \iRF_stage/reg_bank/reg_bank[40] ), .D(
        \iRF_stage/reg_bank/reg_bank[8] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1562 ) );
  MX4X1 \iRF_stage/reg_bank/U1602  ( .A(\iRF_stage/reg_bank/reg_bank[105] ), 
        .B(\iRF_stage/reg_bank/reg_bank[73] ), .C(
        \iRF_stage/reg_bank/reg_bank[41] ), .D(
        \iRF_stage/reg_bank/reg_bank[9] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1572 ) );
  MX4X1 \iRF_stage/reg_bank/U1613  ( .A(\iRF_stage/reg_bank/reg_bank[106] ), 
        .B(\iRF_stage/reg_bank/reg_bank[74] ), .C(
        \iRF_stage/reg_bank/reg_bank[42] ), .D(
        \iRF_stage/reg_bank/reg_bank[10] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1582 ) );
  MX4X1 \iRF_stage/reg_bank/U1624  ( .A(\iRF_stage/reg_bank/reg_bank[107] ), 
        .B(\iRF_stage/reg_bank/reg_bank[75] ), .C(
        \iRF_stage/reg_bank/reg_bank[43] ), .D(
        \iRF_stage/reg_bank/reg_bank[11] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1592 ) );
  MX4X1 \iRF_stage/reg_bank/U1635  ( .A(\iRF_stage/reg_bank/reg_bank[108] ), 
        .B(\iRF_stage/reg_bank/reg_bank[76] ), .C(
        \iRF_stage/reg_bank/reg_bank[44] ), .D(
        \iRF_stage/reg_bank/reg_bank[12] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1602 ) );
  MX4X1 \iRF_stage/reg_bank/U1646  ( .A(\iRF_stage/reg_bank/reg_bank[109] ), 
        .B(\iRF_stage/reg_bank/reg_bank[77] ), .C(
        \iRF_stage/reg_bank/reg_bank[45] ), .D(
        \iRF_stage/reg_bank/reg_bank[13] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1612 ) );
  MX4X1 \iRF_stage/reg_bank/U1657  ( .A(\iRF_stage/reg_bank/reg_bank[110] ), 
        .B(\iRF_stage/reg_bank/reg_bank[78] ), .C(
        \iRF_stage/reg_bank/reg_bank[46] ), .D(
        \iRF_stage/reg_bank/reg_bank[14] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1622 ) );
  MX4X1 \iRF_stage/reg_bank/U1668  ( .A(\iRF_stage/reg_bank/reg_bank[111] ), 
        .B(\iRF_stage/reg_bank/reg_bank[79] ), .C(
        \iRF_stage/reg_bank/reg_bank[47] ), .D(
        \iRF_stage/reg_bank/reg_bank[15] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1632 ) );
  MX4X1 \iRF_stage/reg_bank/U1679  ( .A(\iRF_stage/reg_bank/reg_bank[112] ), 
        .B(\iRF_stage/reg_bank/reg_bank[80] ), .C(
        \iRF_stage/reg_bank/reg_bank[48] ), .D(
        \iRF_stage/reg_bank/reg_bank[16] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1642 ) );
  MX4X1 \iRF_stage/reg_bank/U1690  ( .A(\iRF_stage/reg_bank/reg_bank[113] ), 
        .B(\iRF_stage/reg_bank/reg_bank[81] ), .C(
        \iRF_stage/reg_bank/reg_bank[49] ), .D(
        \iRF_stage/reg_bank/reg_bank[17] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1652 ) );
  MX4X1 \iRF_stage/reg_bank/U1701  ( .A(\iRF_stage/reg_bank/reg_bank[114] ), 
        .B(\iRF_stage/reg_bank/reg_bank[82] ), .C(
        \iRF_stage/reg_bank/reg_bank[50] ), .D(
        \iRF_stage/reg_bank/reg_bank[18] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1662 ) );
  MX4X1 \iRF_stage/reg_bank/U1712  ( .A(\iRF_stage/reg_bank/reg_bank[115] ), 
        .B(\iRF_stage/reg_bank/reg_bank[83] ), .C(
        \iRF_stage/reg_bank/reg_bank[51] ), .D(
        \iRF_stage/reg_bank/reg_bank[19] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1672 ) );
  MX4X1 \iRF_stage/reg_bank/U1723  ( .A(\iRF_stage/reg_bank/reg_bank[116] ), 
        .B(\iRF_stage/reg_bank/reg_bank[84] ), .C(
        \iRF_stage/reg_bank/reg_bank[52] ), .D(
        \iRF_stage/reg_bank/reg_bank[20] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1682 ) );
  MX4X1 \iRF_stage/reg_bank/U1734  ( .A(\iRF_stage/reg_bank/reg_bank[117] ), 
        .B(\iRF_stage/reg_bank/reg_bank[85] ), .C(
        \iRF_stage/reg_bank/reg_bank[53] ), .D(
        \iRF_stage/reg_bank/reg_bank[21] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1692 ) );
  MX4X1 \iRF_stage/reg_bank/U1745  ( .A(\iRF_stage/reg_bank/reg_bank[118] ), 
        .B(\iRF_stage/reg_bank/reg_bank[86] ), .C(
        \iRF_stage/reg_bank/reg_bank[54] ), .D(
        \iRF_stage/reg_bank/reg_bank[22] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1702 ) );
  MX4X1 \iRF_stage/reg_bank/U1756  ( .A(\iRF_stage/reg_bank/reg_bank[119] ), 
        .B(\iRF_stage/reg_bank/reg_bank[87] ), .C(
        \iRF_stage/reg_bank/reg_bank[55] ), .D(
        \iRF_stage/reg_bank/reg_bank[23] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1712 ) );
  MX4X1 \iRF_stage/reg_bank/U1767  ( .A(\iRF_stage/reg_bank/reg_bank[120] ), 
        .B(\iRF_stage/reg_bank/reg_bank[88] ), .C(
        \iRF_stage/reg_bank/reg_bank[56] ), .D(
        \iRF_stage/reg_bank/reg_bank[24] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1722 ) );
  MX4X1 \iRF_stage/reg_bank/U1778  ( .A(\iRF_stage/reg_bank/reg_bank[121] ), 
        .B(\iRF_stage/reg_bank/reg_bank[89] ), .C(
        \iRF_stage/reg_bank/reg_bank[57] ), .D(
        \iRF_stage/reg_bank/reg_bank[25] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1732 ) );
  MX4X1 \iRF_stage/reg_bank/U1789  ( .A(\iRF_stage/reg_bank/reg_bank[122] ), 
        .B(\iRF_stage/reg_bank/reg_bank[90] ), .C(
        \iRF_stage/reg_bank/reg_bank[58] ), .D(
        \iRF_stage/reg_bank/reg_bank[26] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1742 ) );
  MX4X1 \iRF_stage/reg_bank/U1800  ( .A(\iRF_stage/reg_bank/reg_bank[123] ), 
        .B(\iRF_stage/reg_bank/reg_bank[91] ), .C(
        \iRF_stage/reg_bank/reg_bank[59] ), .D(
        \iRF_stage/reg_bank/reg_bank[27] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1752 ) );
  MX4X1 \iRF_stage/reg_bank/U1811  ( .A(\iRF_stage/reg_bank/reg_bank[124] ), 
        .B(\iRF_stage/reg_bank/reg_bank[92] ), .C(
        \iRF_stage/reg_bank/reg_bank[60] ), .D(
        \iRF_stage/reg_bank/reg_bank[28] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1762 ) );
  MX4X1 \iRF_stage/reg_bank/U1822  ( .A(\iRF_stage/reg_bank/reg_bank[125] ), 
        .B(\iRF_stage/reg_bank/reg_bank[93] ), .C(
        \iRF_stage/reg_bank/reg_bank[61] ), .D(
        \iRF_stage/reg_bank/reg_bank[29] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1772 ) );
  MX4X1 \iRF_stage/reg_bank/U1833  ( .A(\iRF_stage/reg_bank/reg_bank[126] ), 
        .B(\iRF_stage/reg_bank/reg_bank[94] ), .C(
        \iRF_stage/reg_bank/reg_bank[62] ), .D(
        \iRF_stage/reg_bank/reg_bank[30] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1782 ) );
  MX4X1 \iRF_stage/reg_bank/U1844  ( .A(\iRF_stage/reg_bank/reg_bank[127] ), 
        .B(\iRF_stage/reg_bank/reg_bank[95] ), .C(
        \iRF_stage/reg_bank/reg_bank[63] ), .D(
        \iRF_stage/reg_bank/reg_bank[31] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1792 ) );
  MX4X1 \iRF_stage/reg_bank/U1151  ( .A(\iRF_stage/reg_bank/reg_bank[96] ), 
        .B(\iRF_stage/reg_bank/reg_bank[64] ), .C(
        \iRF_stage/reg_bank/reg_bank[32] ), .D(
        \iRF_stage/reg_bank/reg_bank[0] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1162 ) );
  MX4X1 \iRF_stage/reg_bank/U1162  ( .A(\iRF_stage/reg_bank/reg_bank[97] ), 
        .B(\iRF_stage/reg_bank/reg_bank[65] ), .C(
        \iRF_stage/reg_bank/reg_bank[33] ), .D(
        \iRF_stage/reg_bank/reg_bank[1] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1172 ) );
  MX4X1 \iRF_stage/reg_bank/U1173  ( .A(\iRF_stage/reg_bank/reg_bank[98] ), 
        .B(\iRF_stage/reg_bank/reg_bank[66] ), .C(
        \iRF_stage/reg_bank/reg_bank[34] ), .D(
        \iRF_stage/reg_bank/reg_bank[2] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1182 ) );
  MX4X1 \iRF_stage/reg_bank/U1184  ( .A(\iRF_stage/reg_bank/reg_bank[99] ), 
        .B(\iRF_stage/reg_bank/reg_bank[67] ), .C(
        \iRF_stage/reg_bank/reg_bank[35] ), .D(
        \iRF_stage/reg_bank/reg_bank[3] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1192 ) );
  MX4X1 \iRF_stage/reg_bank/U1195  ( .A(\iRF_stage/reg_bank/reg_bank[100] ), 
        .B(\iRF_stage/reg_bank/reg_bank[68] ), .C(
        \iRF_stage/reg_bank/reg_bank[36] ), .D(
        \iRF_stage/reg_bank/reg_bank[4] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1202 ) );
  MX4X1 \iRF_stage/reg_bank/U1206  ( .A(\iRF_stage/reg_bank/reg_bank[101] ), 
        .B(\iRF_stage/reg_bank/reg_bank[69] ), .C(
        \iRF_stage/reg_bank/reg_bank[37] ), .D(
        \iRF_stage/reg_bank/reg_bank[5] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1212 ) );
  MX4X1 \iRF_stage/reg_bank/U1217  ( .A(\iRF_stage/reg_bank/reg_bank[102] ), 
        .B(\iRF_stage/reg_bank/reg_bank[70] ), .C(
        \iRF_stage/reg_bank/reg_bank[38] ), .D(
        \iRF_stage/reg_bank/reg_bank[6] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1222 ) );
  MX4X1 \iRF_stage/reg_bank/U1228  ( .A(\iRF_stage/reg_bank/reg_bank[103] ), 
        .B(\iRF_stage/reg_bank/reg_bank[71] ), .C(
        \iRF_stage/reg_bank/reg_bank[39] ), .D(
        \iRF_stage/reg_bank/reg_bank[7] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1232 ) );
  MX4X1 \iRF_stage/reg_bank/U1239  ( .A(\iRF_stage/reg_bank/reg_bank[104] ), 
        .B(\iRF_stage/reg_bank/reg_bank[72] ), .C(
        \iRF_stage/reg_bank/reg_bank[40] ), .D(
        \iRF_stage/reg_bank/reg_bank[8] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1242 ) );
  MX4X1 \iRF_stage/reg_bank/U1250  ( .A(\iRF_stage/reg_bank/reg_bank[105] ), 
        .B(\iRF_stage/reg_bank/reg_bank[73] ), .C(
        \iRF_stage/reg_bank/reg_bank[41] ), .D(
        \iRF_stage/reg_bank/reg_bank[9] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1252 ) );
  MX4X1 \iRF_stage/reg_bank/U1261  ( .A(\iRF_stage/reg_bank/reg_bank[106] ), 
        .B(\iRF_stage/reg_bank/reg_bank[74] ), .C(
        \iRF_stage/reg_bank/reg_bank[42] ), .D(
        \iRF_stage/reg_bank/reg_bank[10] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1262 ) );
  MX4X1 \iRF_stage/reg_bank/U1272  ( .A(\iRF_stage/reg_bank/reg_bank[107] ), 
        .B(\iRF_stage/reg_bank/reg_bank[75] ), .C(
        \iRF_stage/reg_bank/reg_bank[43] ), .D(
        \iRF_stage/reg_bank/reg_bank[11] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1272 ) );
  MX4X1 \iRF_stage/reg_bank/U1283  ( .A(\iRF_stage/reg_bank/reg_bank[108] ), 
        .B(\iRF_stage/reg_bank/reg_bank[76] ), .C(
        \iRF_stage/reg_bank/reg_bank[44] ), .D(
        \iRF_stage/reg_bank/reg_bank[12] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1282 ) );
  MX4X1 \iRF_stage/reg_bank/U1294  ( .A(\iRF_stage/reg_bank/reg_bank[109] ), 
        .B(\iRF_stage/reg_bank/reg_bank[77] ), .C(
        \iRF_stage/reg_bank/reg_bank[45] ), .D(
        \iRF_stage/reg_bank/reg_bank[13] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1292 ) );
  MX4X1 \iRF_stage/reg_bank/U1305  ( .A(\iRF_stage/reg_bank/reg_bank[110] ), 
        .B(\iRF_stage/reg_bank/reg_bank[78] ), .C(
        \iRF_stage/reg_bank/reg_bank[46] ), .D(
        \iRF_stage/reg_bank/reg_bank[14] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1302 ) );
  MX4X1 \iRF_stage/reg_bank/U1316  ( .A(\iRF_stage/reg_bank/reg_bank[111] ), 
        .B(\iRF_stage/reg_bank/reg_bank[79] ), .C(
        \iRF_stage/reg_bank/reg_bank[47] ), .D(
        \iRF_stage/reg_bank/reg_bank[15] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1312 ) );
  MX4X1 \iRF_stage/reg_bank/U1327  ( .A(\iRF_stage/reg_bank/reg_bank[112] ), 
        .B(\iRF_stage/reg_bank/reg_bank[80] ), .C(
        \iRF_stage/reg_bank/reg_bank[48] ), .D(
        \iRF_stage/reg_bank/reg_bank[16] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1322 ) );
  MX4X1 \iRF_stage/reg_bank/U1338  ( .A(\iRF_stage/reg_bank/reg_bank[113] ), 
        .B(\iRF_stage/reg_bank/reg_bank[81] ), .C(
        \iRF_stage/reg_bank/reg_bank[49] ), .D(
        \iRF_stage/reg_bank/reg_bank[17] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1332 ) );
  MX4X1 \iRF_stage/reg_bank/U1349  ( .A(\iRF_stage/reg_bank/reg_bank[114] ), 
        .B(\iRF_stage/reg_bank/reg_bank[82] ), .C(
        \iRF_stage/reg_bank/reg_bank[50] ), .D(
        \iRF_stage/reg_bank/reg_bank[18] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1342 ) );
  MX4X1 \iRF_stage/reg_bank/U1360  ( .A(\iRF_stage/reg_bank/reg_bank[115] ), 
        .B(\iRF_stage/reg_bank/reg_bank[83] ), .C(
        \iRF_stage/reg_bank/reg_bank[51] ), .D(
        \iRF_stage/reg_bank/reg_bank[19] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1352 ) );
  MX4X1 \iRF_stage/reg_bank/U1371  ( .A(\iRF_stage/reg_bank/reg_bank[116] ), 
        .B(\iRF_stage/reg_bank/reg_bank[84] ), .C(
        \iRF_stage/reg_bank/reg_bank[52] ), .D(
        \iRF_stage/reg_bank/reg_bank[20] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1362 ) );
  MX4X1 \iRF_stage/reg_bank/U1382  ( .A(\iRF_stage/reg_bank/reg_bank[117] ), 
        .B(\iRF_stage/reg_bank/reg_bank[85] ), .C(
        \iRF_stage/reg_bank/reg_bank[53] ), .D(
        \iRF_stage/reg_bank/reg_bank[21] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1372 ) );
  MX4X1 \iRF_stage/reg_bank/U1393  ( .A(\iRF_stage/reg_bank/reg_bank[118] ), 
        .B(\iRF_stage/reg_bank/reg_bank[86] ), .C(
        \iRF_stage/reg_bank/reg_bank[54] ), .D(
        \iRF_stage/reg_bank/reg_bank[22] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1382 ) );
  MX4X1 \iRF_stage/reg_bank/U1404  ( .A(\iRF_stage/reg_bank/reg_bank[119] ), 
        .B(\iRF_stage/reg_bank/reg_bank[87] ), .C(
        \iRF_stage/reg_bank/reg_bank[55] ), .D(
        \iRF_stage/reg_bank/reg_bank[23] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1392 ) );
  MX4X1 \iRF_stage/reg_bank/U1415  ( .A(\iRF_stage/reg_bank/reg_bank[120] ), 
        .B(\iRF_stage/reg_bank/reg_bank[88] ), .C(
        \iRF_stage/reg_bank/reg_bank[56] ), .D(
        \iRF_stage/reg_bank/reg_bank[24] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1402 ) );
  MX4X1 \iRF_stage/reg_bank/U1426  ( .A(\iRF_stage/reg_bank/reg_bank[121] ), 
        .B(\iRF_stage/reg_bank/reg_bank[89] ), .C(
        \iRF_stage/reg_bank/reg_bank[57] ), .D(
        \iRF_stage/reg_bank/reg_bank[25] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1412 ) );
  MX4X1 \iRF_stage/reg_bank/U1437  ( .A(\iRF_stage/reg_bank/reg_bank[122] ), 
        .B(\iRF_stage/reg_bank/reg_bank[90] ), .C(
        \iRF_stage/reg_bank/reg_bank[58] ), .D(
        \iRF_stage/reg_bank/reg_bank[26] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1422 ) );
  MX4X1 \iRF_stage/reg_bank/U1448  ( .A(\iRF_stage/reg_bank/reg_bank[123] ), 
        .B(\iRF_stage/reg_bank/reg_bank[91] ), .C(
        \iRF_stage/reg_bank/reg_bank[59] ), .D(
        \iRF_stage/reg_bank/reg_bank[27] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1432 ) );
  MX4X1 \iRF_stage/reg_bank/U1459  ( .A(\iRF_stage/reg_bank/reg_bank[124] ), 
        .B(\iRF_stage/reg_bank/reg_bank[92] ), .C(
        \iRF_stage/reg_bank/reg_bank[60] ), .D(
        \iRF_stage/reg_bank/reg_bank[28] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1442 ) );
  MX4X1 \iRF_stage/reg_bank/U1470  ( .A(\iRF_stage/reg_bank/reg_bank[125] ), 
        .B(\iRF_stage/reg_bank/reg_bank[93] ), .C(
        \iRF_stage/reg_bank/reg_bank[61] ), .D(
        \iRF_stage/reg_bank/reg_bank[29] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1452 ) );
  MX4X1 \iRF_stage/reg_bank/U1481  ( .A(\iRF_stage/reg_bank/reg_bank[126] ), 
        .B(\iRF_stage/reg_bank/reg_bank[94] ), .C(
        \iRF_stage/reg_bank/reg_bank[62] ), .D(
        \iRF_stage/reg_bank/reg_bank[30] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1462 ) );
  MX4X1 \iRF_stage/reg_bank/U1492  ( .A(\iRF_stage/reg_bank/reg_bank[127] ), 
        .B(\iRF_stage/reg_bank/reg_bank[95] ), .C(
        \iRF_stage/reg_bank/reg_bank[63] ), .D(
        \iRF_stage/reg_bank/reg_bank[31] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1472 ) );
  MX4X1 \iRF_stage/reg_bank/U1505  ( .A(\iRF_stage/reg_bank/reg_bank[352] ), 
        .B(\iRF_stage/reg_bank/reg_bank[320] ), .C(
        \iRF_stage/reg_bank/reg_bank[288] ), .D(
        \iRF_stage/reg_bank/reg_bank[256] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1484 ) );
  MX4X1 \iRF_stage/reg_bank/U1510  ( .A(\iRF_stage/reg_bank/reg_bank[864] ), 
        .B(\iRF_stage/reg_bank/reg_bank[832] ), .C(
        \iRF_stage/reg_bank/reg_bank[800] ), .D(
        \iRF_stage/reg_bank/reg_bank[768] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1489 ) );
  MX4X1 \iRF_stage/reg_bank/U1516  ( .A(\iRF_stage/reg_bank/reg_bank[353] ), 
        .B(\iRF_stage/reg_bank/reg_bank[321] ), .C(
        \iRF_stage/reg_bank/reg_bank[289] ), .D(
        \iRF_stage/reg_bank/reg_bank[257] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1494 ) );
  MX4X1 \iRF_stage/reg_bank/U1521  ( .A(\iRF_stage/reg_bank/reg_bank[865] ), 
        .B(\iRF_stage/reg_bank/reg_bank[833] ), .C(
        \iRF_stage/reg_bank/reg_bank[801] ), .D(
        \iRF_stage/reg_bank/reg_bank[769] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1499 ) );
  MX4X1 \iRF_stage/reg_bank/U1527  ( .A(\iRF_stage/reg_bank/reg_bank[354] ), 
        .B(\iRF_stage/reg_bank/reg_bank[322] ), .C(
        \iRF_stage/reg_bank/reg_bank[290] ), .D(
        \iRF_stage/reg_bank/reg_bank[258] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1504 ) );
  MX4X1 \iRF_stage/reg_bank/U1532  ( .A(\iRF_stage/reg_bank/reg_bank[866] ), 
        .B(\iRF_stage/reg_bank/reg_bank[834] ), .C(
        \iRF_stage/reg_bank/reg_bank[802] ), .D(
        \iRF_stage/reg_bank/reg_bank[770] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1509 ) );
  MX4X1 \iRF_stage/reg_bank/U1538  ( .A(\iRF_stage/reg_bank/reg_bank[355] ), 
        .B(\iRF_stage/reg_bank/reg_bank[323] ), .C(
        \iRF_stage/reg_bank/reg_bank[291] ), .D(
        \iRF_stage/reg_bank/reg_bank[259] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1514 ) );
  MX4X1 \iRF_stage/reg_bank/U1543  ( .A(\iRF_stage/reg_bank/reg_bank[867] ), 
        .B(\iRF_stage/reg_bank/reg_bank[835] ), .C(
        \iRF_stage/reg_bank/reg_bank[803] ), .D(
        \iRF_stage/reg_bank/reg_bank[771] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1519 ) );
  MX4X1 \iRF_stage/reg_bank/U1549  ( .A(\iRF_stage/reg_bank/reg_bank[356] ), 
        .B(\iRF_stage/reg_bank/reg_bank[324] ), .C(
        \iRF_stage/reg_bank/reg_bank[292] ), .D(
        \iRF_stage/reg_bank/reg_bank[260] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1524 ) );
  MX4X1 \iRF_stage/reg_bank/U1554  ( .A(\iRF_stage/reg_bank/reg_bank[868] ), 
        .B(\iRF_stage/reg_bank/reg_bank[836] ), .C(
        \iRF_stage/reg_bank/reg_bank[804] ), .D(
        \iRF_stage/reg_bank/reg_bank[772] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1529 ) );
  MX4X1 \iRF_stage/reg_bank/U1560  ( .A(\iRF_stage/reg_bank/reg_bank[357] ), 
        .B(\iRF_stage/reg_bank/reg_bank[325] ), .C(
        \iRF_stage/reg_bank/reg_bank[293] ), .D(
        \iRF_stage/reg_bank/reg_bank[261] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1534 ) );
  MX4X1 \iRF_stage/reg_bank/U1565  ( .A(\iRF_stage/reg_bank/reg_bank[869] ), 
        .B(\iRF_stage/reg_bank/reg_bank[837] ), .C(
        \iRF_stage/reg_bank/reg_bank[805] ), .D(
        \iRF_stage/reg_bank/reg_bank[773] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1539 ) );
  MX4X1 \iRF_stage/reg_bank/U1571  ( .A(\iRF_stage/reg_bank/reg_bank[358] ), 
        .B(\iRF_stage/reg_bank/reg_bank[326] ), .C(
        \iRF_stage/reg_bank/reg_bank[294] ), .D(
        \iRF_stage/reg_bank/reg_bank[262] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1544 ) );
  MX4X1 \iRF_stage/reg_bank/U1576  ( .A(\iRF_stage/reg_bank/reg_bank[870] ), 
        .B(\iRF_stage/reg_bank/reg_bank[838] ), .C(
        \iRF_stage/reg_bank/reg_bank[806] ), .D(
        \iRF_stage/reg_bank/reg_bank[774] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1549 ) );
  MX4X1 \iRF_stage/reg_bank/U1582  ( .A(\iRF_stage/reg_bank/reg_bank[359] ), 
        .B(\iRF_stage/reg_bank/reg_bank[327] ), .C(
        \iRF_stage/reg_bank/reg_bank[295] ), .D(
        \iRF_stage/reg_bank/reg_bank[263] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1554 ) );
  MX4X1 \iRF_stage/reg_bank/U1587  ( .A(\iRF_stage/reg_bank/reg_bank[871] ), 
        .B(\iRF_stage/reg_bank/reg_bank[839] ), .C(
        \iRF_stage/reg_bank/reg_bank[807] ), .D(
        \iRF_stage/reg_bank/reg_bank[775] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1559 ) );
  MX4X1 \iRF_stage/reg_bank/U1593  ( .A(\iRF_stage/reg_bank/reg_bank[360] ), 
        .B(\iRF_stage/reg_bank/reg_bank[328] ), .C(
        \iRF_stage/reg_bank/reg_bank[296] ), .D(
        \iRF_stage/reg_bank/reg_bank[264] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1564 ) );
  MX4X1 \iRF_stage/reg_bank/U1598  ( .A(\iRF_stage/reg_bank/reg_bank[872] ), 
        .B(\iRF_stage/reg_bank/reg_bank[840] ), .C(
        \iRF_stage/reg_bank/reg_bank[808] ), .D(
        \iRF_stage/reg_bank/reg_bank[776] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1569 ) );
  MX4X1 \iRF_stage/reg_bank/U1604  ( .A(\iRF_stage/reg_bank/reg_bank[361] ), 
        .B(\iRF_stage/reg_bank/reg_bank[329] ), .C(
        \iRF_stage/reg_bank/reg_bank[297] ), .D(
        \iRF_stage/reg_bank/reg_bank[265] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1574 ) );
  MX4X1 \iRF_stage/reg_bank/U1609  ( .A(\iRF_stage/reg_bank/reg_bank[873] ), 
        .B(\iRF_stage/reg_bank/reg_bank[841] ), .C(
        \iRF_stage/reg_bank/reg_bank[809] ), .D(
        \iRF_stage/reg_bank/reg_bank[777] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1579 ) );
  MX4X1 \iRF_stage/reg_bank/U1615  ( .A(\iRF_stage/reg_bank/reg_bank[362] ), 
        .B(\iRF_stage/reg_bank/reg_bank[330] ), .C(
        \iRF_stage/reg_bank/reg_bank[298] ), .D(
        \iRF_stage/reg_bank/reg_bank[266] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1584 ) );
  MX4X1 \iRF_stage/reg_bank/U1620  ( .A(\iRF_stage/reg_bank/reg_bank[874] ), 
        .B(\iRF_stage/reg_bank/reg_bank[842] ), .C(
        \iRF_stage/reg_bank/reg_bank[810] ), .D(
        \iRF_stage/reg_bank/reg_bank[778] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1589 ) );
  MX4X1 \iRF_stage/reg_bank/U1626  ( .A(\iRF_stage/reg_bank/reg_bank[363] ), 
        .B(\iRF_stage/reg_bank/reg_bank[331] ), .C(
        \iRF_stage/reg_bank/reg_bank[299] ), .D(
        \iRF_stage/reg_bank/reg_bank[267] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1594 ) );
  MX4X1 \iRF_stage/reg_bank/U1631  ( .A(\iRF_stage/reg_bank/reg_bank[875] ), 
        .B(\iRF_stage/reg_bank/reg_bank[843] ), .C(
        \iRF_stage/reg_bank/reg_bank[811] ), .D(
        \iRF_stage/reg_bank/reg_bank[779] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1599 ) );
  MX4X1 \iRF_stage/reg_bank/U1637  ( .A(\iRF_stage/reg_bank/reg_bank[364] ), 
        .B(\iRF_stage/reg_bank/reg_bank[332] ), .C(
        \iRF_stage/reg_bank/reg_bank[300] ), .D(
        \iRF_stage/reg_bank/reg_bank[268] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1604 ) );
  MX4X1 \iRF_stage/reg_bank/U1642  ( .A(\iRF_stage/reg_bank/reg_bank[876] ), 
        .B(\iRF_stage/reg_bank/reg_bank[844] ), .C(
        \iRF_stage/reg_bank/reg_bank[812] ), .D(
        \iRF_stage/reg_bank/reg_bank[780] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1609 ) );
  MX4X1 \iRF_stage/reg_bank/U1648  ( .A(\iRF_stage/reg_bank/reg_bank[365] ), 
        .B(\iRF_stage/reg_bank/reg_bank[333] ), .C(
        \iRF_stage/reg_bank/reg_bank[301] ), .D(
        \iRF_stage/reg_bank/reg_bank[269] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1614 ) );
  MX4X1 \iRF_stage/reg_bank/U1653  ( .A(\iRF_stage/reg_bank/reg_bank[877] ), 
        .B(\iRF_stage/reg_bank/reg_bank[845] ), .C(
        \iRF_stage/reg_bank/reg_bank[813] ), .D(
        \iRF_stage/reg_bank/reg_bank[781] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1619 ) );
  MX4X1 \iRF_stage/reg_bank/U1659  ( .A(\iRF_stage/reg_bank/reg_bank[366] ), 
        .B(\iRF_stage/reg_bank/reg_bank[334] ), .C(
        \iRF_stage/reg_bank/reg_bank[302] ), .D(
        \iRF_stage/reg_bank/reg_bank[270] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1624 ) );
  MX4X1 \iRF_stage/reg_bank/U1664  ( .A(\iRF_stage/reg_bank/reg_bank[878] ), 
        .B(\iRF_stage/reg_bank/reg_bank[846] ), .C(
        \iRF_stage/reg_bank/reg_bank[814] ), .D(
        \iRF_stage/reg_bank/reg_bank[782] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1629 ) );
  MX4X1 \iRF_stage/reg_bank/U1670  ( .A(\iRF_stage/reg_bank/reg_bank[367] ), 
        .B(\iRF_stage/reg_bank/reg_bank[335] ), .C(
        \iRF_stage/reg_bank/reg_bank[303] ), .D(
        \iRF_stage/reg_bank/reg_bank[271] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1634 ) );
  MX4X1 \iRF_stage/reg_bank/U1675  ( .A(\iRF_stage/reg_bank/reg_bank[879] ), 
        .B(\iRF_stage/reg_bank/reg_bank[847] ), .C(
        \iRF_stage/reg_bank/reg_bank[815] ), .D(
        \iRF_stage/reg_bank/reg_bank[783] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1639 ) );
  MX4X1 \iRF_stage/reg_bank/U1681  ( .A(\iRF_stage/reg_bank/reg_bank[368] ), 
        .B(\iRF_stage/reg_bank/reg_bank[336] ), .C(
        \iRF_stage/reg_bank/reg_bank[304] ), .D(
        \iRF_stage/reg_bank/reg_bank[272] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1644 ) );
  MX4X1 \iRF_stage/reg_bank/U1686  ( .A(\iRF_stage/reg_bank/reg_bank[880] ), 
        .B(\iRF_stage/reg_bank/reg_bank[848] ), .C(
        \iRF_stage/reg_bank/reg_bank[816] ), .D(
        \iRF_stage/reg_bank/reg_bank[784] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1649 ) );
  MX4X1 \iRF_stage/reg_bank/U1692  ( .A(\iRF_stage/reg_bank/reg_bank[369] ), 
        .B(\iRF_stage/reg_bank/reg_bank[337] ), .C(
        \iRF_stage/reg_bank/reg_bank[305] ), .D(
        \iRF_stage/reg_bank/reg_bank[273] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1654 ) );
  MX4X1 \iRF_stage/reg_bank/U1697  ( .A(\iRF_stage/reg_bank/reg_bank[881] ), 
        .B(\iRF_stage/reg_bank/reg_bank[849] ), .C(
        \iRF_stage/reg_bank/reg_bank[817] ), .D(
        \iRF_stage/reg_bank/reg_bank[785] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1659 ) );
  MX4X1 \iRF_stage/reg_bank/U1703  ( .A(\iRF_stage/reg_bank/reg_bank[370] ), 
        .B(\iRF_stage/reg_bank/reg_bank[338] ), .C(
        \iRF_stage/reg_bank/reg_bank[306] ), .D(
        \iRF_stage/reg_bank/reg_bank[274] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1664 ) );
  MX4X1 \iRF_stage/reg_bank/U1708  ( .A(\iRF_stage/reg_bank/reg_bank[882] ), 
        .B(\iRF_stage/reg_bank/reg_bank[850] ), .C(
        \iRF_stage/reg_bank/reg_bank[818] ), .D(
        \iRF_stage/reg_bank/reg_bank[786] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1669 ) );
  MX4X1 \iRF_stage/reg_bank/U1714  ( .A(\iRF_stage/reg_bank/reg_bank[371] ), 
        .B(\iRF_stage/reg_bank/reg_bank[339] ), .C(
        \iRF_stage/reg_bank/reg_bank[307] ), .D(
        \iRF_stage/reg_bank/reg_bank[275] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1674 ) );
  MX4X1 \iRF_stage/reg_bank/U1719  ( .A(\iRF_stage/reg_bank/reg_bank[883] ), 
        .B(\iRF_stage/reg_bank/reg_bank[851] ), .C(
        \iRF_stage/reg_bank/reg_bank[819] ), .D(
        \iRF_stage/reg_bank/reg_bank[787] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1679 ) );
  MX4X1 \iRF_stage/reg_bank/U1725  ( .A(\iRF_stage/reg_bank/reg_bank[372] ), 
        .B(\iRF_stage/reg_bank/reg_bank[340] ), .C(
        \iRF_stage/reg_bank/reg_bank[308] ), .D(
        \iRF_stage/reg_bank/reg_bank[276] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1684 ) );
  MX4X1 \iRF_stage/reg_bank/U1730  ( .A(\iRF_stage/reg_bank/reg_bank[884] ), 
        .B(\iRF_stage/reg_bank/reg_bank[852] ), .C(
        \iRF_stage/reg_bank/reg_bank[820] ), .D(
        \iRF_stage/reg_bank/reg_bank[788] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1689 ) );
  MX4X1 \iRF_stage/reg_bank/U1736  ( .A(\iRF_stage/reg_bank/reg_bank[373] ), 
        .B(\iRF_stage/reg_bank/reg_bank[341] ), .C(
        \iRF_stage/reg_bank/reg_bank[309] ), .D(
        \iRF_stage/reg_bank/reg_bank[277] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1694 ) );
  MX4X1 \iRF_stage/reg_bank/U1741  ( .A(\iRF_stage/reg_bank/reg_bank[885] ), 
        .B(\iRF_stage/reg_bank/reg_bank[853] ), .C(
        \iRF_stage/reg_bank/reg_bank[821] ), .D(
        \iRF_stage/reg_bank/reg_bank[789] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1699 ) );
  MX4X1 \iRF_stage/reg_bank/U1747  ( .A(\iRF_stage/reg_bank/reg_bank[374] ), 
        .B(\iRF_stage/reg_bank/reg_bank[342] ), .C(
        \iRF_stage/reg_bank/reg_bank[310] ), .D(
        \iRF_stage/reg_bank/reg_bank[278] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1704 ) );
  MX4X1 \iRF_stage/reg_bank/U1752  ( .A(\iRF_stage/reg_bank/reg_bank[886] ), 
        .B(\iRF_stage/reg_bank/reg_bank[854] ), .C(
        \iRF_stage/reg_bank/reg_bank[822] ), .D(
        \iRF_stage/reg_bank/reg_bank[790] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1709 ) );
  MX4X1 \iRF_stage/reg_bank/U1758  ( .A(\iRF_stage/reg_bank/reg_bank[375] ), 
        .B(\iRF_stage/reg_bank/reg_bank[343] ), .C(
        \iRF_stage/reg_bank/reg_bank[311] ), .D(
        \iRF_stage/reg_bank/reg_bank[279] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1714 ) );
  MX4X1 \iRF_stage/reg_bank/U1763  ( .A(\iRF_stage/reg_bank/reg_bank[887] ), 
        .B(\iRF_stage/reg_bank/reg_bank[855] ), .C(
        \iRF_stage/reg_bank/reg_bank[823] ), .D(
        \iRF_stage/reg_bank/reg_bank[791] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1719 ) );
  MX4X1 \iRF_stage/reg_bank/U1769  ( .A(\iRF_stage/reg_bank/reg_bank[376] ), 
        .B(\iRF_stage/reg_bank/reg_bank[344] ), .C(
        \iRF_stage/reg_bank/reg_bank[312] ), .D(
        \iRF_stage/reg_bank/reg_bank[280] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1724 ) );
  MX4X1 \iRF_stage/reg_bank/U1774  ( .A(\iRF_stage/reg_bank/reg_bank[888] ), 
        .B(\iRF_stage/reg_bank/reg_bank[856] ), .C(
        \iRF_stage/reg_bank/reg_bank[824] ), .D(
        \iRF_stage/reg_bank/reg_bank[792] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1729 ) );
  MX4X1 \iRF_stage/reg_bank/U1780  ( .A(\iRF_stage/reg_bank/reg_bank[377] ), 
        .B(\iRF_stage/reg_bank/reg_bank[345] ), .C(
        \iRF_stage/reg_bank/reg_bank[313] ), .D(
        \iRF_stage/reg_bank/reg_bank[281] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1734 ) );
  MX4X1 \iRF_stage/reg_bank/U1785  ( .A(\iRF_stage/reg_bank/reg_bank[889] ), 
        .B(\iRF_stage/reg_bank/reg_bank[857] ), .C(
        \iRF_stage/reg_bank/reg_bank[825] ), .D(
        \iRF_stage/reg_bank/reg_bank[793] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1739 ) );
  MX4X1 \iRF_stage/reg_bank/U1791  ( .A(\iRF_stage/reg_bank/reg_bank[378] ), 
        .B(\iRF_stage/reg_bank/reg_bank[346] ), .C(
        \iRF_stage/reg_bank/reg_bank[314] ), .D(
        \iRF_stage/reg_bank/reg_bank[282] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1744 ) );
  MX4X1 \iRF_stage/reg_bank/U1796  ( .A(\iRF_stage/reg_bank/reg_bank[890] ), 
        .B(\iRF_stage/reg_bank/reg_bank[858] ), .C(
        \iRF_stage/reg_bank/reg_bank[826] ), .D(
        \iRF_stage/reg_bank/reg_bank[794] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1749 ) );
  MX4X1 \iRF_stage/reg_bank/U1802  ( .A(\iRF_stage/reg_bank/reg_bank[379] ), 
        .B(\iRF_stage/reg_bank/reg_bank[347] ), .C(
        \iRF_stage/reg_bank/reg_bank[315] ), .D(
        \iRF_stage/reg_bank/reg_bank[283] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1754 ) );
  MX4X1 \iRF_stage/reg_bank/U1807  ( .A(\iRF_stage/reg_bank/reg_bank[891] ), 
        .B(\iRF_stage/reg_bank/reg_bank[859] ), .C(
        \iRF_stage/reg_bank/reg_bank[827] ), .D(
        \iRF_stage/reg_bank/reg_bank[795] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1759 ) );
  MX4X1 \iRF_stage/reg_bank/U1813  ( .A(\iRF_stage/reg_bank/reg_bank[380] ), 
        .B(\iRF_stage/reg_bank/reg_bank[348] ), .C(
        \iRF_stage/reg_bank/reg_bank[316] ), .D(
        \iRF_stage/reg_bank/reg_bank[284] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1764 ) );
  MX4X1 \iRF_stage/reg_bank/U1818  ( .A(\iRF_stage/reg_bank/reg_bank[892] ), 
        .B(\iRF_stage/reg_bank/reg_bank[860] ), .C(
        \iRF_stage/reg_bank/reg_bank[828] ), .D(
        \iRF_stage/reg_bank/reg_bank[796] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1769 ) );
  MX4X1 \iRF_stage/reg_bank/U1824  ( .A(\iRF_stage/reg_bank/reg_bank[381] ), 
        .B(\iRF_stage/reg_bank/reg_bank[349] ), .C(
        \iRF_stage/reg_bank/reg_bank[317] ), .D(
        \iRF_stage/reg_bank/reg_bank[285] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1774 ) );
  MX4X1 \iRF_stage/reg_bank/U1829  ( .A(\iRF_stage/reg_bank/reg_bank[893] ), 
        .B(\iRF_stage/reg_bank/reg_bank[861] ), .C(
        \iRF_stage/reg_bank/reg_bank[829] ), .D(
        \iRF_stage/reg_bank/reg_bank[797] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1779 ) );
  MX4X1 \iRF_stage/reg_bank/U1835  ( .A(\iRF_stage/reg_bank/reg_bank[382] ), 
        .B(\iRF_stage/reg_bank/reg_bank[350] ), .C(
        \iRF_stage/reg_bank/reg_bank[318] ), .D(
        \iRF_stage/reg_bank/reg_bank[286] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1784 ) );
  MX4X1 \iRF_stage/reg_bank/U1840  ( .A(\iRF_stage/reg_bank/reg_bank[894] ), 
        .B(\iRF_stage/reg_bank/reg_bank[862] ), .C(
        \iRF_stage/reg_bank/reg_bank[830] ), .D(
        \iRF_stage/reg_bank/reg_bank[798] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1789 ) );
  MX4X1 \iRF_stage/reg_bank/U1846  ( .A(\iRF_stage/reg_bank/reg_bank[383] ), 
        .B(\iRF_stage/reg_bank/reg_bank[351] ), .C(
        \iRF_stage/reg_bank/reg_bank[319] ), .D(
        \iRF_stage/reg_bank/reg_bank[287] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1794 ) );
  MX4X1 \iRF_stage/reg_bank/U1851  ( .A(\iRF_stage/reg_bank/reg_bank[895] ), 
        .B(\iRF_stage/reg_bank/reg_bank[863] ), .C(
        \iRF_stage/reg_bank/reg_bank[831] ), .D(
        \iRF_stage/reg_bank/reg_bank[799] ), .S0(n247), .S1(
        \iRF_stage/reg_bank/N18 ), .Y(\iRF_stage/reg_bank/n1799 ) );
  MX4X1 \iRF_stage/reg_bank/U1153  ( .A(\iRF_stage/reg_bank/reg_bank[352] ), 
        .B(\iRF_stage/reg_bank/reg_bank[320] ), .C(
        \iRF_stage/reg_bank/reg_bank[288] ), .D(
        \iRF_stage/reg_bank/reg_bank[256] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1164 ) );
  MX4X1 \iRF_stage/reg_bank/U1158  ( .A(\iRF_stage/reg_bank/reg_bank[864] ), 
        .B(\iRF_stage/reg_bank/reg_bank[832] ), .C(
        \iRF_stage/reg_bank/reg_bank[800] ), .D(
        \iRF_stage/reg_bank/reg_bank[768] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1169 ) );
  MX4X1 \iRF_stage/reg_bank/U1164  ( .A(\iRF_stage/reg_bank/reg_bank[353] ), 
        .B(\iRF_stage/reg_bank/reg_bank[321] ), .C(
        \iRF_stage/reg_bank/reg_bank[289] ), .D(
        \iRF_stage/reg_bank/reg_bank[257] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1174 ) );
  MX4X1 \iRF_stage/reg_bank/U1169  ( .A(\iRF_stage/reg_bank/reg_bank[865] ), 
        .B(\iRF_stage/reg_bank/reg_bank[833] ), .C(
        \iRF_stage/reg_bank/reg_bank[801] ), .D(
        \iRF_stage/reg_bank/reg_bank[769] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1179 ) );
  MX4X1 \iRF_stage/reg_bank/U1175  ( .A(\iRF_stage/reg_bank/reg_bank[354] ), 
        .B(\iRF_stage/reg_bank/reg_bank[322] ), .C(
        \iRF_stage/reg_bank/reg_bank[290] ), .D(
        \iRF_stage/reg_bank/reg_bank[258] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1184 ) );
  MX4X1 \iRF_stage/reg_bank/U1180  ( .A(\iRF_stage/reg_bank/reg_bank[866] ), 
        .B(\iRF_stage/reg_bank/reg_bank[834] ), .C(
        \iRF_stage/reg_bank/reg_bank[802] ), .D(
        \iRF_stage/reg_bank/reg_bank[770] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1189 ) );
  MX4X1 \iRF_stage/reg_bank/U1186  ( .A(\iRF_stage/reg_bank/reg_bank[355] ), 
        .B(\iRF_stage/reg_bank/reg_bank[323] ), .C(
        \iRF_stage/reg_bank/reg_bank[291] ), .D(
        \iRF_stage/reg_bank/reg_bank[259] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1194 ) );
  MX4X1 \iRF_stage/reg_bank/U1191  ( .A(\iRF_stage/reg_bank/reg_bank[867] ), 
        .B(\iRF_stage/reg_bank/reg_bank[835] ), .C(
        \iRF_stage/reg_bank/reg_bank[803] ), .D(
        \iRF_stage/reg_bank/reg_bank[771] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1199 ) );
  MX4X1 \iRF_stage/reg_bank/U1197  ( .A(\iRF_stage/reg_bank/reg_bank[356] ), 
        .B(\iRF_stage/reg_bank/reg_bank[324] ), .C(
        \iRF_stage/reg_bank/reg_bank[292] ), .D(
        \iRF_stage/reg_bank/reg_bank[260] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1204 ) );
  MX4X1 \iRF_stage/reg_bank/U1202  ( .A(\iRF_stage/reg_bank/reg_bank[868] ), 
        .B(\iRF_stage/reg_bank/reg_bank[836] ), .C(
        \iRF_stage/reg_bank/reg_bank[804] ), .D(
        \iRF_stage/reg_bank/reg_bank[772] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1209 ) );
  MX4X1 \iRF_stage/reg_bank/U1208  ( .A(\iRF_stage/reg_bank/reg_bank[357] ), 
        .B(\iRF_stage/reg_bank/reg_bank[325] ), .C(
        \iRF_stage/reg_bank/reg_bank[293] ), .D(
        \iRF_stage/reg_bank/reg_bank[261] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1214 ) );
  MX4X1 \iRF_stage/reg_bank/U1213  ( .A(\iRF_stage/reg_bank/reg_bank[869] ), 
        .B(\iRF_stage/reg_bank/reg_bank[837] ), .C(
        \iRF_stage/reg_bank/reg_bank[805] ), .D(
        \iRF_stage/reg_bank/reg_bank[773] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1219 ) );
  MX4X1 \iRF_stage/reg_bank/U1219  ( .A(\iRF_stage/reg_bank/reg_bank[358] ), 
        .B(\iRF_stage/reg_bank/reg_bank[326] ), .C(
        \iRF_stage/reg_bank/reg_bank[294] ), .D(
        \iRF_stage/reg_bank/reg_bank[262] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1224 ) );
  MX4X1 \iRF_stage/reg_bank/U1224  ( .A(\iRF_stage/reg_bank/reg_bank[870] ), 
        .B(\iRF_stage/reg_bank/reg_bank[838] ), .C(
        \iRF_stage/reg_bank/reg_bank[806] ), .D(
        \iRF_stage/reg_bank/reg_bank[774] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1229 ) );
  MX4X1 \iRF_stage/reg_bank/U1230  ( .A(\iRF_stage/reg_bank/reg_bank[359] ), 
        .B(\iRF_stage/reg_bank/reg_bank[327] ), .C(
        \iRF_stage/reg_bank/reg_bank[295] ), .D(
        \iRF_stage/reg_bank/reg_bank[263] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1234 ) );
  MX4X1 \iRF_stage/reg_bank/U1235  ( .A(\iRF_stage/reg_bank/reg_bank[871] ), 
        .B(\iRF_stage/reg_bank/reg_bank[839] ), .C(
        \iRF_stage/reg_bank/reg_bank[807] ), .D(
        \iRF_stage/reg_bank/reg_bank[775] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1239 ) );
  MX4X1 \iRF_stage/reg_bank/U1241  ( .A(\iRF_stage/reg_bank/reg_bank[360] ), 
        .B(\iRF_stage/reg_bank/reg_bank[328] ), .C(
        \iRF_stage/reg_bank/reg_bank[296] ), .D(
        \iRF_stage/reg_bank/reg_bank[264] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1244 ) );
  MX4X1 \iRF_stage/reg_bank/U1246  ( .A(\iRF_stage/reg_bank/reg_bank[872] ), 
        .B(\iRF_stage/reg_bank/reg_bank[840] ), .C(
        \iRF_stage/reg_bank/reg_bank[808] ), .D(
        \iRF_stage/reg_bank/reg_bank[776] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1249 ) );
  MX4X1 \iRF_stage/reg_bank/U1252  ( .A(\iRF_stage/reg_bank/reg_bank[361] ), 
        .B(\iRF_stage/reg_bank/reg_bank[329] ), .C(
        \iRF_stage/reg_bank/reg_bank[297] ), .D(
        \iRF_stage/reg_bank/reg_bank[265] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1254 ) );
  MX4X1 \iRF_stage/reg_bank/U1257  ( .A(\iRF_stage/reg_bank/reg_bank[873] ), 
        .B(\iRF_stage/reg_bank/reg_bank[841] ), .C(
        \iRF_stage/reg_bank/reg_bank[809] ), .D(
        \iRF_stage/reg_bank/reg_bank[777] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1259 ) );
  MX4X1 \iRF_stage/reg_bank/U1263  ( .A(\iRF_stage/reg_bank/reg_bank[362] ), 
        .B(\iRF_stage/reg_bank/reg_bank[330] ), .C(
        \iRF_stage/reg_bank/reg_bank[298] ), .D(
        \iRF_stage/reg_bank/reg_bank[266] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1264 ) );
  MX4X1 \iRF_stage/reg_bank/U1268  ( .A(\iRF_stage/reg_bank/reg_bank[874] ), 
        .B(\iRF_stage/reg_bank/reg_bank[842] ), .C(
        \iRF_stage/reg_bank/reg_bank[810] ), .D(
        \iRF_stage/reg_bank/reg_bank[778] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1269 ) );
  MX4X1 \iRF_stage/reg_bank/U1274  ( .A(\iRF_stage/reg_bank/reg_bank[363] ), 
        .B(\iRF_stage/reg_bank/reg_bank[331] ), .C(
        \iRF_stage/reg_bank/reg_bank[299] ), .D(
        \iRF_stage/reg_bank/reg_bank[267] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1274 ) );
  MX4X1 \iRF_stage/reg_bank/U1279  ( .A(\iRF_stage/reg_bank/reg_bank[875] ), 
        .B(\iRF_stage/reg_bank/reg_bank[843] ), .C(
        \iRF_stage/reg_bank/reg_bank[811] ), .D(
        \iRF_stage/reg_bank/reg_bank[779] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1279 ) );
  MX4X1 \iRF_stage/reg_bank/U1285  ( .A(\iRF_stage/reg_bank/reg_bank[364] ), 
        .B(\iRF_stage/reg_bank/reg_bank[332] ), .C(
        \iRF_stage/reg_bank/reg_bank[300] ), .D(
        \iRF_stage/reg_bank/reg_bank[268] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1284 ) );
  MX4X1 \iRF_stage/reg_bank/U1290  ( .A(\iRF_stage/reg_bank/reg_bank[876] ), 
        .B(\iRF_stage/reg_bank/reg_bank[844] ), .C(
        \iRF_stage/reg_bank/reg_bank[812] ), .D(
        \iRF_stage/reg_bank/reg_bank[780] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1289 ) );
  MX4X1 \iRF_stage/reg_bank/U1296  ( .A(\iRF_stage/reg_bank/reg_bank[365] ), 
        .B(\iRF_stage/reg_bank/reg_bank[333] ), .C(
        \iRF_stage/reg_bank/reg_bank[301] ), .D(
        \iRF_stage/reg_bank/reg_bank[269] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1294 ) );
  MX4X1 \iRF_stage/reg_bank/U1301  ( .A(\iRF_stage/reg_bank/reg_bank[877] ), 
        .B(\iRF_stage/reg_bank/reg_bank[845] ), .C(
        \iRF_stage/reg_bank/reg_bank[813] ), .D(
        \iRF_stage/reg_bank/reg_bank[781] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1299 ) );
  MX4X1 \iRF_stage/reg_bank/U1307  ( .A(\iRF_stage/reg_bank/reg_bank[366] ), 
        .B(\iRF_stage/reg_bank/reg_bank[334] ), .C(
        \iRF_stage/reg_bank/reg_bank[302] ), .D(
        \iRF_stage/reg_bank/reg_bank[270] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1304 ) );
  MX4X1 \iRF_stage/reg_bank/U1312  ( .A(\iRF_stage/reg_bank/reg_bank[878] ), 
        .B(\iRF_stage/reg_bank/reg_bank[846] ), .C(
        \iRF_stage/reg_bank/reg_bank[814] ), .D(
        \iRF_stage/reg_bank/reg_bank[782] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1309 ) );
  MX4X1 \iRF_stage/reg_bank/U1318  ( .A(\iRF_stage/reg_bank/reg_bank[367] ), 
        .B(\iRF_stage/reg_bank/reg_bank[335] ), .C(
        \iRF_stage/reg_bank/reg_bank[303] ), .D(
        \iRF_stage/reg_bank/reg_bank[271] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1314 ) );
  MX4X1 \iRF_stage/reg_bank/U1323  ( .A(\iRF_stage/reg_bank/reg_bank[879] ), 
        .B(\iRF_stage/reg_bank/reg_bank[847] ), .C(
        \iRF_stage/reg_bank/reg_bank[815] ), .D(
        \iRF_stage/reg_bank/reg_bank[783] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1319 ) );
  MX4X1 \iRF_stage/reg_bank/U1329  ( .A(\iRF_stage/reg_bank/reg_bank[368] ), 
        .B(\iRF_stage/reg_bank/reg_bank[336] ), .C(
        \iRF_stage/reg_bank/reg_bank[304] ), .D(
        \iRF_stage/reg_bank/reg_bank[272] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1324 ) );
  MX4X1 \iRF_stage/reg_bank/U1334  ( .A(\iRF_stage/reg_bank/reg_bank[880] ), 
        .B(\iRF_stage/reg_bank/reg_bank[848] ), .C(
        \iRF_stage/reg_bank/reg_bank[816] ), .D(
        \iRF_stage/reg_bank/reg_bank[784] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1329 ) );
  MX4X1 \iRF_stage/reg_bank/U1340  ( .A(\iRF_stage/reg_bank/reg_bank[369] ), 
        .B(\iRF_stage/reg_bank/reg_bank[337] ), .C(
        \iRF_stage/reg_bank/reg_bank[305] ), .D(
        \iRF_stage/reg_bank/reg_bank[273] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1334 ) );
  MX4X1 \iRF_stage/reg_bank/U1345  ( .A(\iRF_stage/reg_bank/reg_bank[881] ), 
        .B(\iRF_stage/reg_bank/reg_bank[849] ), .C(
        \iRF_stage/reg_bank/reg_bank[817] ), .D(
        \iRF_stage/reg_bank/reg_bank[785] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1339 ) );
  MX4X1 \iRF_stage/reg_bank/U1351  ( .A(\iRF_stage/reg_bank/reg_bank[370] ), 
        .B(\iRF_stage/reg_bank/reg_bank[338] ), .C(
        \iRF_stage/reg_bank/reg_bank[306] ), .D(
        \iRF_stage/reg_bank/reg_bank[274] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1344 ) );
  MX4X1 \iRF_stage/reg_bank/U1356  ( .A(\iRF_stage/reg_bank/reg_bank[882] ), 
        .B(\iRF_stage/reg_bank/reg_bank[850] ), .C(
        \iRF_stage/reg_bank/reg_bank[818] ), .D(
        \iRF_stage/reg_bank/reg_bank[786] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1349 ) );
  MX4X1 \iRF_stage/reg_bank/U1362  ( .A(\iRF_stage/reg_bank/reg_bank[371] ), 
        .B(\iRF_stage/reg_bank/reg_bank[339] ), .C(
        \iRF_stage/reg_bank/reg_bank[307] ), .D(
        \iRF_stage/reg_bank/reg_bank[275] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1354 ) );
  MX4X1 \iRF_stage/reg_bank/U1367  ( .A(\iRF_stage/reg_bank/reg_bank[883] ), 
        .B(\iRF_stage/reg_bank/reg_bank[851] ), .C(
        \iRF_stage/reg_bank/reg_bank[819] ), .D(
        \iRF_stage/reg_bank/reg_bank[787] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1359 ) );
  MX4X1 \iRF_stage/reg_bank/U1373  ( .A(\iRF_stage/reg_bank/reg_bank[372] ), 
        .B(\iRF_stage/reg_bank/reg_bank[340] ), .C(
        \iRF_stage/reg_bank/reg_bank[308] ), .D(
        \iRF_stage/reg_bank/reg_bank[276] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1364 ) );
  MX4X1 \iRF_stage/reg_bank/U1378  ( .A(\iRF_stage/reg_bank/reg_bank[884] ), 
        .B(\iRF_stage/reg_bank/reg_bank[852] ), .C(
        \iRF_stage/reg_bank/reg_bank[820] ), .D(
        \iRF_stage/reg_bank/reg_bank[788] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1369 ) );
  MX4X1 \iRF_stage/reg_bank/U1384  ( .A(\iRF_stage/reg_bank/reg_bank[373] ), 
        .B(\iRF_stage/reg_bank/reg_bank[341] ), .C(
        \iRF_stage/reg_bank/reg_bank[309] ), .D(
        \iRF_stage/reg_bank/reg_bank[277] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1374 ) );
  MX4X1 \iRF_stage/reg_bank/U1389  ( .A(\iRF_stage/reg_bank/reg_bank[885] ), 
        .B(\iRF_stage/reg_bank/reg_bank[853] ), .C(
        \iRF_stage/reg_bank/reg_bank[821] ), .D(
        \iRF_stage/reg_bank/reg_bank[789] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1379 ) );
  MX4X1 \iRF_stage/reg_bank/U1395  ( .A(\iRF_stage/reg_bank/reg_bank[374] ), 
        .B(\iRF_stage/reg_bank/reg_bank[342] ), .C(
        \iRF_stage/reg_bank/reg_bank[310] ), .D(
        \iRF_stage/reg_bank/reg_bank[278] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1384 ) );
  MX4X1 \iRF_stage/reg_bank/U1400  ( .A(\iRF_stage/reg_bank/reg_bank[886] ), 
        .B(\iRF_stage/reg_bank/reg_bank[854] ), .C(
        \iRF_stage/reg_bank/reg_bank[822] ), .D(
        \iRF_stage/reg_bank/reg_bank[790] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1389 ) );
  MX4X1 \iRF_stage/reg_bank/U1406  ( .A(\iRF_stage/reg_bank/reg_bank[375] ), 
        .B(\iRF_stage/reg_bank/reg_bank[343] ), .C(
        \iRF_stage/reg_bank/reg_bank[311] ), .D(
        \iRF_stage/reg_bank/reg_bank[279] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1394 ) );
  MX4X1 \iRF_stage/reg_bank/U1411  ( .A(\iRF_stage/reg_bank/reg_bank[887] ), 
        .B(\iRF_stage/reg_bank/reg_bank[855] ), .C(
        \iRF_stage/reg_bank/reg_bank[823] ), .D(
        \iRF_stage/reg_bank/reg_bank[791] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1399 ) );
  MX4X1 \iRF_stage/reg_bank/U1417  ( .A(\iRF_stage/reg_bank/reg_bank[376] ), 
        .B(\iRF_stage/reg_bank/reg_bank[344] ), .C(
        \iRF_stage/reg_bank/reg_bank[312] ), .D(
        \iRF_stage/reg_bank/reg_bank[280] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1404 ) );
  MX4X1 \iRF_stage/reg_bank/U1422  ( .A(\iRF_stage/reg_bank/reg_bank[888] ), 
        .B(\iRF_stage/reg_bank/reg_bank[856] ), .C(
        \iRF_stage/reg_bank/reg_bank[824] ), .D(
        \iRF_stage/reg_bank/reg_bank[792] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1409 ) );
  MX4X1 \iRF_stage/reg_bank/U1428  ( .A(\iRF_stage/reg_bank/reg_bank[377] ), 
        .B(\iRF_stage/reg_bank/reg_bank[345] ), .C(
        \iRF_stage/reg_bank/reg_bank[313] ), .D(
        \iRF_stage/reg_bank/reg_bank[281] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1414 ) );
  MX4X1 \iRF_stage/reg_bank/U1433  ( .A(\iRF_stage/reg_bank/reg_bank[889] ), 
        .B(\iRF_stage/reg_bank/reg_bank[857] ), .C(
        \iRF_stage/reg_bank/reg_bank[825] ), .D(
        \iRF_stage/reg_bank/reg_bank[793] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1419 ) );
  MX4X1 \iRF_stage/reg_bank/U1439  ( .A(\iRF_stage/reg_bank/reg_bank[378] ), 
        .B(\iRF_stage/reg_bank/reg_bank[346] ), .C(
        \iRF_stage/reg_bank/reg_bank[314] ), .D(
        \iRF_stage/reg_bank/reg_bank[282] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1424 ) );
  MX4X1 \iRF_stage/reg_bank/U1444  ( .A(\iRF_stage/reg_bank/reg_bank[890] ), 
        .B(\iRF_stage/reg_bank/reg_bank[858] ), .C(
        \iRF_stage/reg_bank/reg_bank[826] ), .D(
        \iRF_stage/reg_bank/reg_bank[794] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1429 ) );
  MX4X1 \iRF_stage/reg_bank/U1450  ( .A(\iRF_stage/reg_bank/reg_bank[379] ), 
        .B(\iRF_stage/reg_bank/reg_bank[347] ), .C(
        \iRF_stage/reg_bank/reg_bank[315] ), .D(
        \iRF_stage/reg_bank/reg_bank[283] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1434 ) );
  MX4X1 \iRF_stage/reg_bank/U1455  ( .A(\iRF_stage/reg_bank/reg_bank[891] ), 
        .B(\iRF_stage/reg_bank/reg_bank[859] ), .C(
        \iRF_stage/reg_bank/reg_bank[827] ), .D(
        \iRF_stage/reg_bank/reg_bank[795] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1439 ) );
  MX4X1 \iRF_stage/reg_bank/U1461  ( .A(\iRF_stage/reg_bank/reg_bank[380] ), 
        .B(\iRF_stage/reg_bank/reg_bank[348] ), .C(
        \iRF_stage/reg_bank/reg_bank[316] ), .D(
        \iRF_stage/reg_bank/reg_bank[284] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1444 ) );
  MX4X1 \iRF_stage/reg_bank/U1466  ( .A(\iRF_stage/reg_bank/reg_bank[892] ), 
        .B(\iRF_stage/reg_bank/reg_bank[860] ), .C(
        \iRF_stage/reg_bank/reg_bank[828] ), .D(
        \iRF_stage/reg_bank/reg_bank[796] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1449 ) );
  MX4X1 \iRF_stage/reg_bank/U1472  ( .A(\iRF_stage/reg_bank/reg_bank[381] ), 
        .B(\iRF_stage/reg_bank/reg_bank[349] ), .C(
        \iRF_stage/reg_bank/reg_bank[317] ), .D(
        \iRF_stage/reg_bank/reg_bank[285] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1454 ) );
  MX4X1 \iRF_stage/reg_bank/U1477  ( .A(\iRF_stage/reg_bank/reg_bank[893] ), 
        .B(\iRF_stage/reg_bank/reg_bank[861] ), .C(
        \iRF_stage/reg_bank/reg_bank[829] ), .D(
        \iRF_stage/reg_bank/reg_bank[797] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1459 ) );
  MX4X1 \iRF_stage/reg_bank/U1483  ( .A(\iRF_stage/reg_bank/reg_bank[382] ), 
        .B(\iRF_stage/reg_bank/reg_bank[350] ), .C(
        \iRF_stage/reg_bank/reg_bank[318] ), .D(
        \iRF_stage/reg_bank/reg_bank[286] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1464 ) );
  MX4X1 \iRF_stage/reg_bank/U1488  ( .A(\iRF_stage/reg_bank/reg_bank[894] ), 
        .B(\iRF_stage/reg_bank/reg_bank[862] ), .C(
        \iRF_stage/reg_bank/reg_bank[830] ), .D(
        \iRF_stage/reg_bank/reg_bank[798] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1469 ) );
  MX4X1 \iRF_stage/reg_bank/U1494  ( .A(\iRF_stage/reg_bank/reg_bank[383] ), 
        .B(\iRF_stage/reg_bank/reg_bank[351] ), .C(
        \iRF_stage/reg_bank/reg_bank[319] ), .D(
        \iRF_stage/reg_bank/reg_bank[287] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1474 ) );
  MX4X1 \iRF_stage/reg_bank/U1499  ( .A(\iRF_stage/reg_bank/reg_bank[895] ), 
        .B(\iRF_stage/reg_bank/reg_bank[863] ), .C(
        \iRF_stage/reg_bank/reg_bank[831] ), .D(
        \iRF_stage/reg_bank/reg_bank[799] ), .S0(n197), .S1(
        \iRF_stage/reg_bank/N13 ), .Y(\iRF_stage/reg_bank/n1479 ) );
  MX4X1 \iRF_stage/reg_bank/U1508  ( .A(\iRF_stage/reg_bank/reg_bank[608] ), 
        .B(\iRF_stage/reg_bank/reg_bank[576] ), .C(
        \iRF_stage/reg_bank/reg_bank[544] ), .D(
        \iRF_stage/reg_bank/reg_bank[512] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1487 ) );
  MX4X1 \iRF_stage/reg_bank/U1511  ( .A(\iRF_stage/reg_bank/reg_bank[992] ), 
        .B(\iRF_stage/reg_bank/reg_bank[960] ), .C(
        \iRF_stage/reg_bank/reg_bank[928] ), .D(
        \iRF_stage/reg_bank/reg_bank[896] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1490 ) );
  MX4X1 \iRF_stage/reg_bank/U1509  ( .A(\iRF_stage/reg_bank/reg_bank[736] ), 
        .B(\iRF_stage/reg_bank/reg_bank[704] ), .C(
        \iRF_stage/reg_bank/reg_bank[672] ), .D(
        \iRF_stage/reg_bank/reg_bank[640] ), .S0(n226), .S1(n251), .Y(
        \iRF_stage/reg_bank/n1488 ) );
  MX4XL \iRF_stage/reg_bank/U1512  ( .A(\iRF_stage/reg_bank/n1490 ), .B(
        \iRF_stage/reg_bank/n1488 ), .C(\iRF_stage/reg_bank/n1489 ), .D(
        \iRF_stage/reg_bank/n1487 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1491 ) );
  MX4X1 \iRF_stage/reg_bank/U1519  ( .A(\iRF_stage/reg_bank/reg_bank[609] ), 
        .B(\iRF_stage/reg_bank/reg_bank[577] ), .C(
        \iRF_stage/reg_bank/reg_bank[545] ), .D(
        \iRF_stage/reg_bank/reg_bank[513] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1497 ) );
  MX4X1 \iRF_stage/reg_bank/U1522  ( .A(\iRF_stage/reg_bank/reg_bank[993] ), 
        .B(\iRF_stage/reg_bank/reg_bank[961] ), .C(
        \iRF_stage/reg_bank/reg_bank[929] ), .D(
        \iRF_stage/reg_bank/reg_bank[897] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1500 ) );
  MX4X1 \iRF_stage/reg_bank/U1520  ( .A(\iRF_stage/reg_bank/reg_bank[737] ), 
        .B(\iRF_stage/reg_bank/reg_bank[705] ), .C(
        \iRF_stage/reg_bank/reg_bank[673] ), .D(
        \iRF_stage/reg_bank/reg_bank[641] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1498 ) );
  MX4XL \iRF_stage/reg_bank/U1523  ( .A(\iRF_stage/reg_bank/n1500 ), .B(
        \iRF_stage/reg_bank/n1498 ), .C(\iRF_stage/reg_bank/n1499 ), .D(
        \iRF_stage/reg_bank/n1497 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1501 ) );
  MX4X1 \iRF_stage/reg_bank/U1530  ( .A(\iRF_stage/reg_bank/reg_bank[610] ), 
        .B(\iRF_stage/reg_bank/reg_bank[578] ), .C(
        \iRF_stage/reg_bank/reg_bank[546] ), .D(
        \iRF_stage/reg_bank/reg_bank[514] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1507 ) );
  MX4X1 \iRF_stage/reg_bank/U1533  ( .A(\iRF_stage/reg_bank/reg_bank[994] ), 
        .B(\iRF_stage/reg_bank/reg_bank[962] ), .C(
        \iRF_stage/reg_bank/reg_bank[930] ), .D(
        \iRF_stage/reg_bank/reg_bank[898] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1510 ) );
  MX4X1 \iRF_stage/reg_bank/U1531  ( .A(\iRF_stage/reg_bank/reg_bank[738] ), 
        .B(\iRF_stage/reg_bank/reg_bank[706] ), .C(
        \iRF_stage/reg_bank/reg_bank[674] ), .D(
        \iRF_stage/reg_bank/reg_bank[642] ), .S0(n227), .S1(n252), .Y(
        \iRF_stage/reg_bank/n1508 ) );
  MX4XL \iRF_stage/reg_bank/U1534  ( .A(\iRF_stage/reg_bank/n1510 ), .B(
        \iRF_stage/reg_bank/n1508 ), .C(\iRF_stage/reg_bank/n1509 ), .D(
        \iRF_stage/reg_bank/n1507 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1511 ) );
  MX4X1 \iRF_stage/reg_bank/U1541  ( .A(\iRF_stage/reg_bank/reg_bank[611] ), 
        .B(\iRF_stage/reg_bank/reg_bank[579] ), .C(
        \iRF_stage/reg_bank/reg_bank[547] ), .D(
        \iRF_stage/reg_bank/reg_bank[515] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1517 ) );
  MX4X1 \iRF_stage/reg_bank/U1544  ( .A(\iRF_stage/reg_bank/reg_bank[995] ), 
        .B(\iRF_stage/reg_bank/reg_bank[963] ), .C(
        \iRF_stage/reg_bank/reg_bank[931] ), .D(
        \iRF_stage/reg_bank/reg_bank[899] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1520 ) );
  MX4X1 \iRF_stage/reg_bank/U1542  ( .A(\iRF_stage/reg_bank/reg_bank[739] ), 
        .B(\iRF_stage/reg_bank/reg_bank[707] ), .C(
        \iRF_stage/reg_bank/reg_bank[675] ), .D(
        \iRF_stage/reg_bank/reg_bank[643] ), .S0(n228), .S1(n253), .Y(
        \iRF_stage/reg_bank/n1518 ) );
  MX4XL \iRF_stage/reg_bank/U1545  ( .A(\iRF_stage/reg_bank/n1520 ), .B(
        \iRF_stage/reg_bank/n1518 ), .C(\iRF_stage/reg_bank/n1519 ), .D(
        \iRF_stage/reg_bank/n1517 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1521 ) );
  MX4X1 \iRF_stage/reg_bank/U1552  ( .A(\iRF_stage/reg_bank/reg_bank[612] ), 
        .B(\iRF_stage/reg_bank/reg_bank[580] ), .C(
        \iRF_stage/reg_bank/reg_bank[548] ), .D(
        \iRF_stage/reg_bank/reg_bank[516] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1527 ) );
  MX4X1 \iRF_stage/reg_bank/U1555  ( .A(\iRF_stage/reg_bank/reg_bank[996] ), 
        .B(\iRF_stage/reg_bank/reg_bank[964] ), .C(
        \iRF_stage/reg_bank/reg_bank[932] ), .D(
        \iRF_stage/reg_bank/reg_bank[900] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1530 ) );
  MX4X1 \iRF_stage/reg_bank/U1553  ( .A(\iRF_stage/reg_bank/reg_bank[740] ), 
        .B(\iRF_stage/reg_bank/reg_bank[708] ), .C(
        \iRF_stage/reg_bank/reg_bank[676] ), .D(
        \iRF_stage/reg_bank/reg_bank[644] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1528 ) );
  MX4XL \iRF_stage/reg_bank/U1556  ( .A(\iRF_stage/reg_bank/n1530 ), .B(
        \iRF_stage/reg_bank/n1528 ), .C(\iRF_stage/reg_bank/n1529 ), .D(
        \iRF_stage/reg_bank/n1527 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1531 ) );
  MX4X1 \iRF_stage/reg_bank/U1563  ( .A(\iRF_stage/reg_bank/reg_bank[613] ), 
        .B(\iRF_stage/reg_bank/reg_bank[581] ), .C(
        \iRF_stage/reg_bank/reg_bank[549] ), .D(
        \iRF_stage/reg_bank/reg_bank[517] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1537 ) );
  MX4X1 \iRF_stage/reg_bank/U1566  ( .A(\iRF_stage/reg_bank/reg_bank[997] ), 
        .B(\iRF_stage/reg_bank/reg_bank[965] ), .C(
        \iRF_stage/reg_bank/reg_bank[933] ), .D(
        \iRF_stage/reg_bank/reg_bank[901] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1540 ) );
  MX4X1 \iRF_stage/reg_bank/U1564  ( .A(\iRF_stage/reg_bank/reg_bank[741] ), 
        .B(\iRF_stage/reg_bank/reg_bank[709] ), .C(
        \iRF_stage/reg_bank/reg_bank[677] ), .D(
        \iRF_stage/reg_bank/reg_bank[645] ), .S0(n229), .S1(n254), .Y(
        \iRF_stage/reg_bank/n1538 ) );
  MX4XL \iRF_stage/reg_bank/U1567  ( .A(\iRF_stage/reg_bank/n1540 ), .B(
        \iRF_stage/reg_bank/n1538 ), .C(\iRF_stage/reg_bank/n1539 ), .D(
        \iRF_stage/reg_bank/n1537 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1541 ) );
  MX4X1 \iRF_stage/reg_bank/U1574  ( .A(\iRF_stage/reg_bank/reg_bank[614] ), 
        .B(\iRF_stage/reg_bank/reg_bank[582] ), .C(
        \iRF_stage/reg_bank/reg_bank[550] ), .D(
        \iRF_stage/reg_bank/reg_bank[518] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1547 ) );
  MX4X1 \iRF_stage/reg_bank/U1577  ( .A(\iRF_stage/reg_bank/reg_bank[998] ), 
        .B(\iRF_stage/reg_bank/reg_bank[966] ), .C(
        \iRF_stage/reg_bank/reg_bank[934] ), .D(
        \iRF_stage/reg_bank/reg_bank[902] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1550 ) );
  MX4X1 \iRF_stage/reg_bank/U1575  ( .A(\iRF_stage/reg_bank/reg_bank[742] ), 
        .B(\iRF_stage/reg_bank/reg_bank[710] ), .C(
        \iRF_stage/reg_bank/reg_bank[678] ), .D(
        \iRF_stage/reg_bank/reg_bank[646] ), .S0(n230), .S1(n255), .Y(
        \iRF_stage/reg_bank/n1548 ) );
  MX4XL \iRF_stage/reg_bank/U1578  ( .A(\iRF_stage/reg_bank/n1550 ), .B(
        \iRF_stage/reg_bank/n1548 ), .C(\iRF_stage/reg_bank/n1549 ), .D(
        \iRF_stage/reg_bank/n1547 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1551 ) );
  MX4X1 \iRF_stage/reg_bank/U1585  ( .A(\iRF_stage/reg_bank/reg_bank[615] ), 
        .B(\iRF_stage/reg_bank/reg_bank[583] ), .C(
        \iRF_stage/reg_bank/reg_bank[551] ), .D(
        \iRF_stage/reg_bank/reg_bank[519] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1557 ) );
  MX4X1 \iRF_stage/reg_bank/U1588  ( .A(\iRF_stage/reg_bank/reg_bank[999] ), 
        .B(\iRF_stage/reg_bank/reg_bank[967] ), .C(
        \iRF_stage/reg_bank/reg_bank[935] ), .D(
        \iRF_stage/reg_bank/reg_bank[903] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1560 ) );
  MX4X1 \iRF_stage/reg_bank/U1586  ( .A(\iRF_stage/reg_bank/reg_bank[743] ), 
        .B(\iRF_stage/reg_bank/reg_bank[711] ), .C(
        \iRF_stage/reg_bank/reg_bank[679] ), .D(
        \iRF_stage/reg_bank/reg_bank[647] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1558 ) );
  MX4XL \iRF_stage/reg_bank/U1589  ( .A(\iRF_stage/reg_bank/n1560 ), .B(
        \iRF_stage/reg_bank/n1558 ), .C(\iRF_stage/reg_bank/n1559 ), .D(
        \iRF_stage/reg_bank/n1557 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1561 ) );
  MX4X1 \iRF_stage/reg_bank/U1596  ( .A(\iRF_stage/reg_bank/reg_bank[616] ), 
        .B(\iRF_stage/reg_bank/reg_bank[584] ), .C(
        \iRF_stage/reg_bank/reg_bank[552] ), .D(
        \iRF_stage/reg_bank/reg_bank[520] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1567 ) );
  MX4X1 \iRF_stage/reg_bank/U1599  ( .A(\iRF_stage/reg_bank/reg_bank[1000] ), 
        .B(\iRF_stage/reg_bank/reg_bank[968] ), .C(
        \iRF_stage/reg_bank/reg_bank[936] ), .D(
        \iRF_stage/reg_bank/reg_bank[904] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1570 ) );
  MX4X1 \iRF_stage/reg_bank/U1597  ( .A(\iRF_stage/reg_bank/reg_bank[744] ), 
        .B(\iRF_stage/reg_bank/reg_bank[712] ), .C(
        \iRF_stage/reg_bank/reg_bank[680] ), .D(
        \iRF_stage/reg_bank/reg_bank[648] ), .S0(n231), .S1(n256), .Y(
        \iRF_stage/reg_bank/n1568 ) );
  MX4XL \iRF_stage/reg_bank/U1600  ( .A(\iRF_stage/reg_bank/n1570 ), .B(
        \iRF_stage/reg_bank/n1568 ), .C(\iRF_stage/reg_bank/n1569 ), .D(
        \iRF_stage/reg_bank/n1567 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1571 ) );
  MX4X1 \iRF_stage/reg_bank/U1607  ( .A(\iRF_stage/reg_bank/reg_bank[617] ), 
        .B(\iRF_stage/reg_bank/reg_bank[585] ), .C(
        \iRF_stage/reg_bank/reg_bank[553] ), .D(
        \iRF_stage/reg_bank/reg_bank[521] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1577 ) );
  MX4X1 \iRF_stage/reg_bank/U1610  ( .A(\iRF_stage/reg_bank/reg_bank[1001] ), 
        .B(\iRF_stage/reg_bank/reg_bank[969] ), .C(
        \iRF_stage/reg_bank/reg_bank[937] ), .D(
        \iRF_stage/reg_bank/reg_bank[905] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1580 ) );
  MX4X1 \iRF_stage/reg_bank/U1608  ( .A(\iRF_stage/reg_bank/reg_bank[745] ), 
        .B(\iRF_stage/reg_bank/reg_bank[713] ), .C(
        \iRF_stage/reg_bank/reg_bank[681] ), .D(
        \iRF_stage/reg_bank/reg_bank[649] ), .S0(n232), .S1(n257), .Y(
        \iRF_stage/reg_bank/n1578 ) );
  MX4XL \iRF_stage/reg_bank/U1611  ( .A(\iRF_stage/reg_bank/n1580 ), .B(
        \iRF_stage/reg_bank/n1578 ), .C(\iRF_stage/reg_bank/n1579 ), .D(
        \iRF_stage/reg_bank/n1577 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1581 ) );
  MX4X1 \iRF_stage/reg_bank/U1618  ( .A(\iRF_stage/reg_bank/reg_bank[618] ), 
        .B(\iRF_stage/reg_bank/reg_bank[586] ), .C(
        \iRF_stage/reg_bank/reg_bank[554] ), .D(
        \iRF_stage/reg_bank/reg_bank[522] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1587 ) );
  MX4X1 \iRF_stage/reg_bank/U1621  ( .A(\iRF_stage/reg_bank/reg_bank[1002] ), 
        .B(\iRF_stage/reg_bank/reg_bank[970] ), .C(
        \iRF_stage/reg_bank/reg_bank[938] ), .D(
        \iRF_stage/reg_bank/reg_bank[906] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1590 ) );
  MX4X1 \iRF_stage/reg_bank/U1619  ( .A(\iRF_stage/reg_bank/reg_bank[746] ), 
        .B(\iRF_stage/reg_bank/reg_bank[714] ), .C(
        \iRF_stage/reg_bank/reg_bank[682] ), .D(
        \iRF_stage/reg_bank/reg_bank[650] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1588 ) );
  MX4XL \iRF_stage/reg_bank/U1622  ( .A(\iRF_stage/reg_bank/n1590 ), .B(
        \iRF_stage/reg_bank/n1588 ), .C(\iRF_stage/reg_bank/n1589 ), .D(
        \iRF_stage/reg_bank/n1587 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1591 ) );
  MX4X1 \iRF_stage/reg_bank/U1629  ( .A(\iRF_stage/reg_bank/reg_bank[619] ), 
        .B(\iRF_stage/reg_bank/reg_bank[587] ), .C(
        \iRF_stage/reg_bank/reg_bank[555] ), .D(
        \iRF_stage/reg_bank/reg_bank[523] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1597 ) );
  MX4X1 \iRF_stage/reg_bank/U1632  ( .A(\iRF_stage/reg_bank/reg_bank[1003] ), 
        .B(\iRF_stage/reg_bank/reg_bank[971] ), .C(
        \iRF_stage/reg_bank/reg_bank[939] ), .D(
        \iRF_stage/reg_bank/reg_bank[907] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1600 ) );
  MX4X1 \iRF_stage/reg_bank/U1630  ( .A(\iRF_stage/reg_bank/reg_bank[747] ), 
        .B(\iRF_stage/reg_bank/reg_bank[715] ), .C(
        \iRF_stage/reg_bank/reg_bank[683] ), .D(
        \iRF_stage/reg_bank/reg_bank[651] ), .S0(n233), .S1(n258), .Y(
        \iRF_stage/reg_bank/n1598 ) );
  MX4XL \iRF_stage/reg_bank/U1633  ( .A(\iRF_stage/reg_bank/n1600 ), .B(
        \iRF_stage/reg_bank/n1598 ), .C(\iRF_stage/reg_bank/n1599 ), .D(
        \iRF_stage/reg_bank/n1597 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1601 ) );
  MX4X1 \iRF_stage/reg_bank/U1640  ( .A(\iRF_stage/reg_bank/reg_bank[620] ), 
        .B(\iRF_stage/reg_bank/reg_bank[588] ), .C(
        \iRF_stage/reg_bank/reg_bank[556] ), .D(
        \iRF_stage/reg_bank/reg_bank[524] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1607 ) );
  MX4X1 \iRF_stage/reg_bank/U1643  ( .A(\iRF_stage/reg_bank/reg_bank[1004] ), 
        .B(\iRF_stage/reg_bank/reg_bank[972] ), .C(
        \iRF_stage/reg_bank/reg_bank[940] ), .D(
        \iRF_stage/reg_bank/reg_bank[908] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1610 ) );
  MX4X1 \iRF_stage/reg_bank/U1641  ( .A(\iRF_stage/reg_bank/reg_bank[748] ), 
        .B(\iRF_stage/reg_bank/reg_bank[716] ), .C(
        \iRF_stage/reg_bank/reg_bank[684] ), .D(
        \iRF_stage/reg_bank/reg_bank[652] ), .S0(n234), .S1(n259), .Y(
        \iRF_stage/reg_bank/n1608 ) );
  MX4XL \iRF_stage/reg_bank/U1644  ( .A(\iRF_stage/reg_bank/n1610 ), .B(
        \iRF_stage/reg_bank/n1608 ), .C(\iRF_stage/reg_bank/n1609 ), .D(
        \iRF_stage/reg_bank/n1607 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1611 ) );
  MX4X1 \iRF_stage/reg_bank/U1651  ( .A(\iRF_stage/reg_bank/reg_bank[621] ), 
        .B(\iRF_stage/reg_bank/reg_bank[589] ), .C(
        \iRF_stage/reg_bank/reg_bank[557] ), .D(
        \iRF_stage/reg_bank/reg_bank[525] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1617 ) );
  MX4X1 \iRF_stage/reg_bank/U1654  ( .A(\iRF_stage/reg_bank/reg_bank[1005] ), 
        .B(\iRF_stage/reg_bank/reg_bank[973] ), .C(
        \iRF_stage/reg_bank/reg_bank[941] ), .D(
        \iRF_stage/reg_bank/reg_bank[909] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1620 ) );
  MX4X1 \iRF_stage/reg_bank/U1652  ( .A(\iRF_stage/reg_bank/reg_bank[749] ), 
        .B(\iRF_stage/reg_bank/reg_bank[717] ), .C(
        \iRF_stage/reg_bank/reg_bank[685] ), .D(
        \iRF_stage/reg_bank/reg_bank[653] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1618 ) );
  MX4XL \iRF_stage/reg_bank/U1655  ( .A(\iRF_stage/reg_bank/n1620 ), .B(
        \iRF_stage/reg_bank/n1618 ), .C(\iRF_stage/reg_bank/n1619 ), .D(
        \iRF_stage/reg_bank/n1617 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1621 ) );
  MX4X1 \iRF_stage/reg_bank/U1662  ( .A(\iRF_stage/reg_bank/reg_bank[622] ), 
        .B(\iRF_stage/reg_bank/reg_bank[590] ), .C(
        \iRF_stage/reg_bank/reg_bank[558] ), .D(
        \iRF_stage/reg_bank/reg_bank[526] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1627 ) );
  MX4X1 \iRF_stage/reg_bank/U1665  ( .A(\iRF_stage/reg_bank/reg_bank[1006] ), 
        .B(\iRF_stage/reg_bank/reg_bank[974] ), .C(
        \iRF_stage/reg_bank/reg_bank[942] ), .D(
        \iRF_stage/reg_bank/reg_bank[910] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1630 ) );
  MX4X1 \iRF_stage/reg_bank/U1663  ( .A(\iRF_stage/reg_bank/reg_bank[750] ), 
        .B(\iRF_stage/reg_bank/reg_bank[718] ), .C(
        \iRF_stage/reg_bank/reg_bank[686] ), .D(
        \iRF_stage/reg_bank/reg_bank[654] ), .S0(n235), .S1(n260), .Y(
        \iRF_stage/reg_bank/n1628 ) );
  MX4XL \iRF_stage/reg_bank/U1666  ( .A(\iRF_stage/reg_bank/n1630 ), .B(
        \iRF_stage/reg_bank/n1628 ), .C(\iRF_stage/reg_bank/n1629 ), .D(
        \iRF_stage/reg_bank/n1627 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1631 ) );
  MX4X1 \iRF_stage/reg_bank/U1673  ( .A(\iRF_stage/reg_bank/reg_bank[623] ), 
        .B(\iRF_stage/reg_bank/reg_bank[591] ), .C(
        \iRF_stage/reg_bank/reg_bank[559] ), .D(
        \iRF_stage/reg_bank/reg_bank[527] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1637 ) );
  MX4X1 \iRF_stage/reg_bank/U1676  ( .A(\iRF_stage/reg_bank/reg_bank[1007] ), 
        .B(\iRF_stage/reg_bank/reg_bank[975] ), .C(
        \iRF_stage/reg_bank/reg_bank[943] ), .D(
        \iRF_stage/reg_bank/reg_bank[911] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1640 ) );
  MX4X1 \iRF_stage/reg_bank/U1674  ( .A(\iRF_stage/reg_bank/reg_bank[751] ), 
        .B(\iRF_stage/reg_bank/reg_bank[719] ), .C(
        \iRF_stage/reg_bank/reg_bank[687] ), .D(
        \iRF_stage/reg_bank/reg_bank[655] ), .S0(n236), .S1(n261), .Y(
        \iRF_stage/reg_bank/n1638 ) );
  MX4XL \iRF_stage/reg_bank/U1677  ( .A(\iRF_stage/reg_bank/n1640 ), .B(
        \iRF_stage/reg_bank/n1638 ), .C(\iRF_stage/reg_bank/n1639 ), .D(
        \iRF_stage/reg_bank/n1637 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1641 ) );
  MX4X1 \iRF_stage/reg_bank/U1684  ( .A(\iRF_stage/reg_bank/reg_bank[624] ), 
        .B(\iRF_stage/reg_bank/reg_bank[592] ), .C(
        \iRF_stage/reg_bank/reg_bank[560] ), .D(
        \iRF_stage/reg_bank/reg_bank[528] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1647 ) );
  MX4X1 \iRF_stage/reg_bank/U1687  ( .A(\iRF_stage/reg_bank/reg_bank[1008] ), 
        .B(\iRF_stage/reg_bank/reg_bank[976] ), .C(
        \iRF_stage/reg_bank/reg_bank[944] ), .D(
        \iRF_stage/reg_bank/reg_bank[912] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1650 ) );
  MX4X1 \iRF_stage/reg_bank/U1685  ( .A(\iRF_stage/reg_bank/reg_bank[752] ), 
        .B(\iRF_stage/reg_bank/reg_bank[720] ), .C(
        \iRF_stage/reg_bank/reg_bank[688] ), .D(
        \iRF_stage/reg_bank/reg_bank[656] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1648 ) );
  MX4XL \iRF_stage/reg_bank/U1688  ( .A(\iRF_stage/reg_bank/n1650 ), .B(
        \iRF_stage/reg_bank/n1648 ), .C(\iRF_stage/reg_bank/n1649 ), .D(
        \iRF_stage/reg_bank/n1647 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1651 ) );
  MX4X1 \iRF_stage/reg_bank/U1695  ( .A(\iRF_stage/reg_bank/reg_bank[625] ), 
        .B(\iRF_stage/reg_bank/reg_bank[593] ), .C(
        \iRF_stage/reg_bank/reg_bank[561] ), .D(
        \iRF_stage/reg_bank/reg_bank[529] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1657 ) );
  MX4X1 \iRF_stage/reg_bank/U1698  ( .A(\iRF_stage/reg_bank/reg_bank[1009] ), 
        .B(\iRF_stage/reg_bank/reg_bank[977] ), .C(
        \iRF_stage/reg_bank/reg_bank[945] ), .D(
        \iRF_stage/reg_bank/reg_bank[913] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1660 ) );
  MX4X1 \iRF_stage/reg_bank/U1696  ( .A(\iRF_stage/reg_bank/reg_bank[753] ), 
        .B(\iRF_stage/reg_bank/reg_bank[721] ), .C(
        \iRF_stage/reg_bank/reg_bank[689] ), .D(
        \iRF_stage/reg_bank/reg_bank[657] ), .S0(n237), .S1(n262), .Y(
        \iRF_stage/reg_bank/n1658 ) );
  MX4XL \iRF_stage/reg_bank/U1699  ( .A(\iRF_stage/reg_bank/n1660 ), .B(
        \iRF_stage/reg_bank/n1658 ), .C(\iRF_stage/reg_bank/n1659 ), .D(
        \iRF_stage/reg_bank/n1657 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1661 ) );
  MX4X1 \iRF_stage/reg_bank/U1706  ( .A(\iRF_stage/reg_bank/reg_bank[626] ), 
        .B(\iRF_stage/reg_bank/reg_bank[594] ), .C(
        \iRF_stage/reg_bank/reg_bank[562] ), .D(
        \iRF_stage/reg_bank/reg_bank[530] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1667 ) );
  MX4X1 \iRF_stage/reg_bank/U1709  ( .A(\iRF_stage/reg_bank/reg_bank[1010] ), 
        .B(\iRF_stage/reg_bank/reg_bank[978] ), .C(
        \iRF_stage/reg_bank/reg_bank[946] ), .D(
        \iRF_stage/reg_bank/reg_bank[914] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1670 ) );
  MX4X1 \iRF_stage/reg_bank/U1707  ( .A(\iRF_stage/reg_bank/reg_bank[754] ), 
        .B(\iRF_stage/reg_bank/reg_bank[722] ), .C(
        \iRF_stage/reg_bank/reg_bank[690] ), .D(
        \iRF_stage/reg_bank/reg_bank[658] ), .S0(n238), .S1(n263), .Y(
        \iRF_stage/reg_bank/n1668 ) );
  MX4XL \iRF_stage/reg_bank/U1710  ( .A(\iRF_stage/reg_bank/n1670 ), .B(
        \iRF_stage/reg_bank/n1668 ), .C(\iRF_stage/reg_bank/n1669 ), .D(
        \iRF_stage/reg_bank/n1667 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1671 ) );
  MX4X1 \iRF_stage/reg_bank/U1717  ( .A(\iRF_stage/reg_bank/reg_bank[627] ), 
        .B(\iRF_stage/reg_bank/reg_bank[595] ), .C(
        \iRF_stage/reg_bank/reg_bank[563] ), .D(
        \iRF_stage/reg_bank/reg_bank[531] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1677 ) );
  MX4X1 \iRF_stage/reg_bank/U1720  ( .A(\iRF_stage/reg_bank/reg_bank[1011] ), 
        .B(\iRF_stage/reg_bank/reg_bank[979] ), .C(
        \iRF_stage/reg_bank/reg_bank[947] ), .D(
        \iRF_stage/reg_bank/reg_bank[915] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1680 ) );
  MX4X1 \iRF_stage/reg_bank/U1718  ( .A(\iRF_stage/reg_bank/reg_bank[755] ), 
        .B(\iRF_stage/reg_bank/reg_bank[723] ), .C(
        \iRF_stage/reg_bank/reg_bank[691] ), .D(
        \iRF_stage/reg_bank/reg_bank[659] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1678 ) );
  MX4XL \iRF_stage/reg_bank/U1721  ( .A(\iRF_stage/reg_bank/n1680 ), .B(
        \iRF_stage/reg_bank/n1678 ), .C(\iRF_stage/reg_bank/n1679 ), .D(
        \iRF_stage/reg_bank/n1677 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1681 ) );
  MX4X1 \iRF_stage/reg_bank/U1728  ( .A(\iRF_stage/reg_bank/reg_bank[628] ), 
        .B(\iRF_stage/reg_bank/reg_bank[596] ), .C(
        \iRF_stage/reg_bank/reg_bank[564] ), .D(
        \iRF_stage/reg_bank/reg_bank[532] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1687 ) );
  MX4X1 \iRF_stage/reg_bank/U1731  ( .A(\iRF_stage/reg_bank/reg_bank[1012] ), 
        .B(\iRF_stage/reg_bank/reg_bank[980] ), .C(
        \iRF_stage/reg_bank/reg_bank[948] ), .D(
        \iRF_stage/reg_bank/reg_bank[916] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1690 ) );
  MX4X1 \iRF_stage/reg_bank/U1729  ( .A(\iRF_stage/reg_bank/reg_bank[756] ), 
        .B(\iRF_stage/reg_bank/reg_bank[724] ), .C(
        \iRF_stage/reg_bank/reg_bank[692] ), .D(
        \iRF_stage/reg_bank/reg_bank[660] ), .S0(n239), .S1(n264), .Y(
        \iRF_stage/reg_bank/n1688 ) );
  MX4XL \iRF_stage/reg_bank/U1732  ( .A(\iRF_stage/reg_bank/n1690 ), .B(
        \iRF_stage/reg_bank/n1688 ), .C(\iRF_stage/reg_bank/n1689 ), .D(
        \iRF_stage/reg_bank/n1687 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1691 ) );
  MX4X1 \iRF_stage/reg_bank/U1739  ( .A(\iRF_stage/reg_bank/reg_bank[629] ), 
        .B(\iRF_stage/reg_bank/reg_bank[597] ), .C(
        \iRF_stage/reg_bank/reg_bank[565] ), .D(
        \iRF_stage/reg_bank/reg_bank[533] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1697 ) );
  MX4X1 \iRF_stage/reg_bank/U1742  ( .A(\iRF_stage/reg_bank/reg_bank[1013] ), 
        .B(\iRF_stage/reg_bank/reg_bank[981] ), .C(
        \iRF_stage/reg_bank/reg_bank[949] ), .D(
        \iRF_stage/reg_bank/reg_bank[917] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1700 ) );
  MX4X1 \iRF_stage/reg_bank/U1740  ( .A(\iRF_stage/reg_bank/reg_bank[757] ), 
        .B(\iRF_stage/reg_bank/reg_bank[725] ), .C(
        \iRF_stage/reg_bank/reg_bank[693] ), .D(
        \iRF_stage/reg_bank/reg_bank[661] ), .S0(n240), .S1(n265), .Y(
        \iRF_stage/reg_bank/n1698 ) );
  MX4XL \iRF_stage/reg_bank/U1743  ( .A(\iRF_stage/reg_bank/n1700 ), .B(
        \iRF_stage/reg_bank/n1698 ), .C(\iRF_stage/reg_bank/n1699 ), .D(
        \iRF_stage/reg_bank/n1697 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1701 ) );
  MX4X1 \iRF_stage/reg_bank/U1750  ( .A(\iRF_stage/reg_bank/reg_bank[630] ), 
        .B(\iRF_stage/reg_bank/reg_bank[598] ), .C(
        \iRF_stage/reg_bank/reg_bank[566] ), .D(
        \iRF_stage/reg_bank/reg_bank[534] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1707 ) );
  MX4X1 \iRF_stage/reg_bank/U1753  ( .A(\iRF_stage/reg_bank/reg_bank[1014] ), 
        .B(\iRF_stage/reg_bank/reg_bank[982] ), .C(
        \iRF_stage/reg_bank/reg_bank[950] ), .D(
        \iRF_stage/reg_bank/reg_bank[918] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1710 ) );
  MX4X1 \iRF_stage/reg_bank/U1751  ( .A(\iRF_stage/reg_bank/reg_bank[758] ), 
        .B(\iRF_stage/reg_bank/reg_bank[726] ), .C(
        \iRF_stage/reg_bank/reg_bank[694] ), .D(
        \iRF_stage/reg_bank/reg_bank[662] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1708 ) );
  MX4XL \iRF_stage/reg_bank/U1754  ( .A(\iRF_stage/reg_bank/n1710 ), .B(
        \iRF_stage/reg_bank/n1708 ), .C(\iRF_stage/reg_bank/n1709 ), .D(
        \iRF_stage/reg_bank/n1707 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1711 ) );
  MX4X1 \iRF_stage/reg_bank/U1761  ( .A(\iRF_stage/reg_bank/reg_bank[631] ), 
        .B(\iRF_stage/reg_bank/reg_bank[599] ), .C(
        \iRF_stage/reg_bank/reg_bank[567] ), .D(
        \iRF_stage/reg_bank/reg_bank[535] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1717 ) );
  MX4X1 \iRF_stage/reg_bank/U1764  ( .A(\iRF_stage/reg_bank/reg_bank[1015] ), 
        .B(\iRF_stage/reg_bank/reg_bank[983] ), .C(
        \iRF_stage/reg_bank/reg_bank[951] ), .D(
        \iRF_stage/reg_bank/reg_bank[919] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1720 ) );
  MX4X1 \iRF_stage/reg_bank/U1762  ( .A(\iRF_stage/reg_bank/reg_bank[759] ), 
        .B(\iRF_stage/reg_bank/reg_bank[727] ), .C(
        \iRF_stage/reg_bank/reg_bank[695] ), .D(
        \iRF_stage/reg_bank/reg_bank[663] ), .S0(n241), .S1(n266), .Y(
        \iRF_stage/reg_bank/n1718 ) );
  MX4XL \iRF_stage/reg_bank/U1765  ( .A(\iRF_stage/reg_bank/n1720 ), .B(
        \iRF_stage/reg_bank/n1718 ), .C(\iRF_stage/reg_bank/n1719 ), .D(
        \iRF_stage/reg_bank/n1717 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1721 ) );
  MX4X1 \iRF_stage/reg_bank/U1772  ( .A(\iRF_stage/reg_bank/reg_bank[632] ), 
        .B(\iRF_stage/reg_bank/reg_bank[600] ), .C(
        \iRF_stage/reg_bank/reg_bank[568] ), .D(
        \iRF_stage/reg_bank/reg_bank[536] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1727 ) );
  MX4X1 \iRF_stage/reg_bank/U1775  ( .A(\iRF_stage/reg_bank/reg_bank[1016] ), 
        .B(\iRF_stage/reg_bank/reg_bank[984] ), .C(
        \iRF_stage/reg_bank/reg_bank[952] ), .D(
        \iRF_stage/reg_bank/reg_bank[920] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1730 ) );
  MX4X1 \iRF_stage/reg_bank/U1773  ( .A(\iRF_stage/reg_bank/reg_bank[760] ), 
        .B(\iRF_stage/reg_bank/reg_bank[728] ), .C(
        \iRF_stage/reg_bank/reg_bank[696] ), .D(
        \iRF_stage/reg_bank/reg_bank[664] ), .S0(n242), .S1(n267), .Y(
        \iRF_stage/reg_bank/n1728 ) );
  MX4XL \iRF_stage/reg_bank/U1776  ( .A(\iRF_stage/reg_bank/n1730 ), .B(
        \iRF_stage/reg_bank/n1728 ), .C(\iRF_stage/reg_bank/n1729 ), .D(
        \iRF_stage/reg_bank/n1727 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1731 ) );
  MX4X1 \iRF_stage/reg_bank/U1783  ( .A(\iRF_stage/reg_bank/reg_bank[633] ), 
        .B(\iRF_stage/reg_bank/reg_bank[601] ), .C(
        \iRF_stage/reg_bank/reg_bank[569] ), .D(
        \iRF_stage/reg_bank/reg_bank[537] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1737 ) );
  MX4X1 \iRF_stage/reg_bank/U1786  ( .A(\iRF_stage/reg_bank/reg_bank[1017] ), 
        .B(\iRF_stage/reg_bank/reg_bank[985] ), .C(
        \iRF_stage/reg_bank/reg_bank[953] ), .D(
        \iRF_stage/reg_bank/reg_bank[921] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1740 ) );
  MX4X1 \iRF_stage/reg_bank/U1784  ( .A(\iRF_stage/reg_bank/reg_bank[761] ), 
        .B(\iRF_stage/reg_bank/reg_bank[729] ), .C(
        \iRF_stage/reg_bank/reg_bank[697] ), .D(
        \iRF_stage/reg_bank/reg_bank[665] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1738 ) );
  MX4XL \iRF_stage/reg_bank/U1787  ( .A(\iRF_stage/reg_bank/n1740 ), .B(
        \iRF_stage/reg_bank/n1738 ), .C(\iRF_stage/reg_bank/n1739 ), .D(
        \iRF_stage/reg_bank/n1737 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1741 ) );
  MX4X1 \iRF_stage/reg_bank/U1794  ( .A(\iRF_stage/reg_bank/reg_bank[634] ), 
        .B(\iRF_stage/reg_bank/reg_bank[602] ), .C(
        \iRF_stage/reg_bank/reg_bank[570] ), .D(
        \iRF_stage/reg_bank/reg_bank[538] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1747 ) );
  MX4X1 \iRF_stage/reg_bank/U1797  ( .A(\iRF_stage/reg_bank/reg_bank[1018] ), 
        .B(\iRF_stage/reg_bank/reg_bank[986] ), .C(
        \iRF_stage/reg_bank/reg_bank[954] ), .D(
        \iRF_stage/reg_bank/reg_bank[922] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1750 ) );
  MX4X1 \iRF_stage/reg_bank/U1795  ( .A(\iRF_stage/reg_bank/reg_bank[762] ), 
        .B(\iRF_stage/reg_bank/reg_bank[730] ), .C(
        \iRF_stage/reg_bank/reg_bank[698] ), .D(
        \iRF_stage/reg_bank/reg_bank[666] ), .S0(n243), .S1(n268), .Y(
        \iRF_stage/reg_bank/n1748 ) );
  MX4XL \iRF_stage/reg_bank/U1798  ( .A(\iRF_stage/reg_bank/n1750 ), .B(
        \iRF_stage/reg_bank/n1748 ), .C(\iRF_stage/reg_bank/n1749 ), .D(
        \iRF_stage/reg_bank/n1747 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1751 ) );
  MX4X1 \iRF_stage/reg_bank/U1805  ( .A(\iRF_stage/reg_bank/reg_bank[635] ), 
        .B(\iRF_stage/reg_bank/reg_bank[603] ), .C(
        \iRF_stage/reg_bank/reg_bank[571] ), .D(
        \iRF_stage/reg_bank/reg_bank[539] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1757 ) );
  MX4X1 \iRF_stage/reg_bank/U1808  ( .A(\iRF_stage/reg_bank/reg_bank[1019] ), 
        .B(\iRF_stage/reg_bank/reg_bank[987] ), .C(
        \iRF_stage/reg_bank/reg_bank[955] ), .D(
        \iRF_stage/reg_bank/reg_bank[923] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1760 ) );
  MX4X1 \iRF_stage/reg_bank/U1806  ( .A(\iRF_stage/reg_bank/reg_bank[763] ), 
        .B(\iRF_stage/reg_bank/reg_bank[731] ), .C(
        \iRF_stage/reg_bank/reg_bank[699] ), .D(
        \iRF_stage/reg_bank/reg_bank[667] ), .S0(n244), .S1(n269), .Y(
        \iRF_stage/reg_bank/n1758 ) );
  MX4XL \iRF_stage/reg_bank/U1809  ( .A(\iRF_stage/reg_bank/n1760 ), .B(
        \iRF_stage/reg_bank/n1758 ), .C(\iRF_stage/reg_bank/n1759 ), .D(
        \iRF_stage/reg_bank/n1757 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1761 ) );
  MX4X1 \iRF_stage/reg_bank/U1816  ( .A(\iRF_stage/reg_bank/reg_bank[636] ), 
        .B(\iRF_stage/reg_bank/reg_bank[604] ), .C(
        \iRF_stage/reg_bank/reg_bank[572] ), .D(
        \iRF_stage/reg_bank/reg_bank[540] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1767 ) );
  MX4X1 \iRF_stage/reg_bank/U1819  ( .A(\iRF_stage/reg_bank/reg_bank[1020] ), 
        .B(\iRF_stage/reg_bank/reg_bank[988] ), .C(
        \iRF_stage/reg_bank/reg_bank[956] ), .D(
        \iRF_stage/reg_bank/reg_bank[924] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1770 ) );
  MX4X1 \iRF_stage/reg_bank/U1817  ( .A(\iRF_stage/reg_bank/reg_bank[764] ), 
        .B(\iRF_stage/reg_bank/reg_bank[732] ), .C(
        \iRF_stage/reg_bank/reg_bank[700] ), .D(
        \iRF_stage/reg_bank/reg_bank[668] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1768 ) );
  MX4XL \iRF_stage/reg_bank/U1820  ( .A(\iRF_stage/reg_bank/n1770 ), .B(
        \iRF_stage/reg_bank/n1768 ), .C(\iRF_stage/reg_bank/n1769 ), .D(
        \iRF_stage/reg_bank/n1767 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1771 ) );
  MX4X1 \iRF_stage/reg_bank/U1827  ( .A(\iRF_stage/reg_bank/reg_bank[637] ), 
        .B(\iRF_stage/reg_bank/reg_bank[605] ), .C(
        \iRF_stage/reg_bank/reg_bank[573] ), .D(
        \iRF_stage/reg_bank/reg_bank[541] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1777 ) );
  MX4X1 \iRF_stage/reg_bank/U1830  ( .A(\iRF_stage/reg_bank/reg_bank[1021] ), 
        .B(\iRF_stage/reg_bank/reg_bank[989] ), .C(
        \iRF_stage/reg_bank/reg_bank[957] ), .D(
        \iRF_stage/reg_bank/reg_bank[925] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1780 ) );
  MX4X1 \iRF_stage/reg_bank/U1828  ( .A(\iRF_stage/reg_bank/reg_bank[765] ), 
        .B(\iRF_stage/reg_bank/reg_bank[733] ), .C(
        \iRF_stage/reg_bank/reg_bank[701] ), .D(
        \iRF_stage/reg_bank/reg_bank[669] ), .S0(n245), .S1(n270), .Y(
        \iRF_stage/reg_bank/n1778 ) );
  MX4XL \iRF_stage/reg_bank/U1831  ( .A(\iRF_stage/reg_bank/n1780 ), .B(
        \iRF_stage/reg_bank/n1778 ), .C(\iRF_stage/reg_bank/n1779 ), .D(
        \iRF_stage/reg_bank/n1777 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1781 ) );
  MX4X1 \iRF_stage/reg_bank/U1838  ( .A(\iRF_stage/reg_bank/reg_bank[638] ), 
        .B(\iRF_stage/reg_bank/reg_bank[606] ), .C(
        \iRF_stage/reg_bank/reg_bank[574] ), .D(
        \iRF_stage/reg_bank/reg_bank[542] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1787 ) );
  MX4X1 \iRF_stage/reg_bank/U1841  ( .A(\iRF_stage/reg_bank/reg_bank[1022] ), 
        .B(\iRF_stage/reg_bank/reg_bank[990] ), .C(
        \iRF_stage/reg_bank/reg_bank[958] ), .D(
        \iRF_stage/reg_bank/reg_bank[926] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1790 ) );
  MX4X1 \iRF_stage/reg_bank/U1839  ( .A(\iRF_stage/reg_bank/reg_bank[766] ), 
        .B(\iRF_stage/reg_bank/reg_bank[734] ), .C(
        \iRF_stage/reg_bank/reg_bank[702] ), .D(
        \iRF_stage/reg_bank/reg_bank[670] ), .S0(n246), .S1(n271), .Y(
        \iRF_stage/reg_bank/n1788 ) );
  MX4XL \iRF_stage/reg_bank/U1842  ( .A(\iRF_stage/reg_bank/n1790 ), .B(
        \iRF_stage/reg_bank/n1788 ), .C(\iRF_stage/reg_bank/n1789 ), .D(
        \iRF_stage/reg_bank/n1787 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1791 ) );
  MX4X1 \iRF_stage/reg_bank/U1849  ( .A(\iRF_stage/reg_bank/reg_bank[639] ), 
        .B(\iRF_stage/reg_bank/reg_bank[607] ), .C(
        \iRF_stage/reg_bank/reg_bank[575] ), .D(
        \iRF_stage/reg_bank/reg_bank[543] ), .S0(n247), .S1(
        \iRF_stage/reg_bank/N18 ), .Y(\iRF_stage/reg_bank/n1797 ) );
  MX4X1 \iRF_stage/reg_bank/U1852  ( .A(\iRF_stage/reg_bank/reg_bank[1023] ), 
        .B(\iRF_stage/reg_bank/reg_bank[991] ), .C(
        \iRF_stage/reg_bank/reg_bank[959] ), .D(
        \iRF_stage/reg_bank/reg_bank[927] ), .S0(n247), .S1(
        \iRF_stage/reg_bank/N18 ), .Y(\iRF_stage/reg_bank/n1800 ) );
  MX4X1 \iRF_stage/reg_bank/U1850  ( .A(\iRF_stage/reg_bank/reg_bank[767] ), 
        .B(\iRF_stage/reg_bank/reg_bank[735] ), .C(
        \iRF_stage/reg_bank/reg_bank[703] ), .D(
        \iRF_stage/reg_bank/reg_bank[671] ), .S0(n247), .S1(
        \iRF_stage/reg_bank/N18 ), .Y(\iRF_stage/reg_bank/n1798 ) );
  MX4X1 \iRF_stage/reg_bank/U1853  ( .A(\iRF_stage/reg_bank/n1800 ), .B(
        \iRF_stage/reg_bank/n1798 ), .C(\iRF_stage/reg_bank/n1799 ), .D(
        \iRF_stage/reg_bank/n1797 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1801 ) );
  MX4X1 \iRF_stage/reg_bank/U1156  ( .A(\iRF_stage/reg_bank/reg_bank[608] ), 
        .B(\iRF_stage/reg_bank/reg_bank[576] ), .C(
        \iRF_stage/reg_bank/reg_bank[544] ), .D(
        \iRF_stage/reg_bank/reg_bank[512] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1167 ) );
  MX4X1 \iRF_stage/reg_bank/U1159  ( .A(\iRF_stage/reg_bank/reg_bank[992] ), 
        .B(\iRF_stage/reg_bank/reg_bank[960] ), .C(
        \iRF_stage/reg_bank/reg_bank[928] ), .D(
        \iRF_stage/reg_bank/reg_bank[896] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1170 ) );
  MX4X1 \iRF_stage/reg_bank/U1157  ( .A(\iRF_stage/reg_bank/reg_bank[736] ), 
        .B(\iRF_stage/reg_bank/reg_bank[704] ), .C(
        \iRF_stage/reg_bank/reg_bank[672] ), .D(
        \iRF_stage/reg_bank/reg_bank[640] ), .S0(n176), .S1(n201), .Y(
        \iRF_stage/reg_bank/n1168 ) );
  MX4XL \iRF_stage/reg_bank/U1160  ( .A(\iRF_stage/reg_bank/n1170 ), .B(
        \iRF_stage/reg_bank/n1168 ), .C(\iRF_stage/reg_bank/n1169 ), .D(
        \iRF_stage/reg_bank/n1167 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1171 ) );
  MX4X1 \iRF_stage/reg_bank/U1167  ( .A(\iRF_stage/reg_bank/reg_bank[609] ), 
        .B(\iRF_stage/reg_bank/reg_bank[577] ), .C(
        \iRF_stage/reg_bank/reg_bank[545] ), .D(
        \iRF_stage/reg_bank/reg_bank[513] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1177 ) );
  MX4X1 \iRF_stage/reg_bank/U1170  ( .A(\iRF_stage/reg_bank/reg_bank[993] ), 
        .B(\iRF_stage/reg_bank/reg_bank[961] ), .C(
        \iRF_stage/reg_bank/reg_bank[929] ), .D(
        \iRF_stage/reg_bank/reg_bank[897] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1180 ) );
  MX4X1 \iRF_stage/reg_bank/U1168  ( .A(\iRF_stage/reg_bank/reg_bank[737] ), 
        .B(\iRF_stage/reg_bank/reg_bank[705] ), .C(
        \iRF_stage/reg_bank/reg_bank[673] ), .D(
        \iRF_stage/reg_bank/reg_bank[641] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1178 ) );
  MX4XL \iRF_stage/reg_bank/U1171  ( .A(\iRF_stage/reg_bank/n1180 ), .B(
        \iRF_stage/reg_bank/n1178 ), .C(\iRF_stage/reg_bank/n1179 ), .D(
        \iRF_stage/reg_bank/n1177 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1181 ) );
  MX4X1 \iRF_stage/reg_bank/U1178  ( .A(\iRF_stage/reg_bank/reg_bank[610] ), 
        .B(\iRF_stage/reg_bank/reg_bank[578] ), .C(
        \iRF_stage/reg_bank/reg_bank[546] ), .D(
        \iRF_stage/reg_bank/reg_bank[514] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1187 ) );
  MX4X1 \iRF_stage/reg_bank/U1181  ( .A(\iRF_stage/reg_bank/reg_bank[994] ), 
        .B(\iRF_stage/reg_bank/reg_bank[962] ), .C(
        \iRF_stage/reg_bank/reg_bank[930] ), .D(
        \iRF_stage/reg_bank/reg_bank[898] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1190 ) );
  MX4X1 \iRF_stage/reg_bank/U1179  ( .A(\iRF_stage/reg_bank/reg_bank[738] ), 
        .B(\iRF_stage/reg_bank/reg_bank[706] ), .C(
        \iRF_stage/reg_bank/reg_bank[674] ), .D(
        \iRF_stage/reg_bank/reg_bank[642] ), .S0(n177), .S1(n202), .Y(
        \iRF_stage/reg_bank/n1188 ) );
  MX4XL \iRF_stage/reg_bank/U1182  ( .A(\iRF_stage/reg_bank/n1190 ), .B(
        \iRF_stage/reg_bank/n1188 ), .C(\iRF_stage/reg_bank/n1189 ), .D(
        \iRF_stage/reg_bank/n1187 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1191 ) );
  MX4X1 \iRF_stage/reg_bank/U1189  ( .A(\iRF_stage/reg_bank/reg_bank[611] ), 
        .B(\iRF_stage/reg_bank/reg_bank[579] ), .C(
        \iRF_stage/reg_bank/reg_bank[547] ), .D(
        \iRF_stage/reg_bank/reg_bank[515] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1197 ) );
  MX4X1 \iRF_stage/reg_bank/U1192  ( .A(\iRF_stage/reg_bank/reg_bank[995] ), 
        .B(\iRF_stage/reg_bank/reg_bank[963] ), .C(
        \iRF_stage/reg_bank/reg_bank[931] ), .D(
        \iRF_stage/reg_bank/reg_bank[899] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1200 ) );
  MX4X1 \iRF_stage/reg_bank/U1190  ( .A(\iRF_stage/reg_bank/reg_bank[739] ), 
        .B(\iRF_stage/reg_bank/reg_bank[707] ), .C(
        \iRF_stage/reg_bank/reg_bank[675] ), .D(
        \iRF_stage/reg_bank/reg_bank[643] ), .S0(n178), .S1(n203), .Y(
        \iRF_stage/reg_bank/n1198 ) );
  MX4XL \iRF_stage/reg_bank/U1193  ( .A(\iRF_stage/reg_bank/n1200 ), .B(
        \iRF_stage/reg_bank/n1198 ), .C(\iRF_stage/reg_bank/n1199 ), .D(
        \iRF_stage/reg_bank/n1197 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1201 ) );
  MX4X1 \iRF_stage/reg_bank/U1200  ( .A(\iRF_stage/reg_bank/reg_bank[612] ), 
        .B(\iRF_stage/reg_bank/reg_bank[580] ), .C(
        \iRF_stage/reg_bank/reg_bank[548] ), .D(
        \iRF_stage/reg_bank/reg_bank[516] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1207 ) );
  MX4X1 \iRF_stage/reg_bank/U1203  ( .A(\iRF_stage/reg_bank/reg_bank[996] ), 
        .B(\iRF_stage/reg_bank/reg_bank[964] ), .C(
        \iRF_stage/reg_bank/reg_bank[932] ), .D(
        \iRF_stage/reg_bank/reg_bank[900] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1210 ) );
  MX4X1 \iRF_stage/reg_bank/U1201  ( .A(\iRF_stage/reg_bank/reg_bank[740] ), 
        .B(\iRF_stage/reg_bank/reg_bank[708] ), .C(
        \iRF_stage/reg_bank/reg_bank[676] ), .D(
        \iRF_stage/reg_bank/reg_bank[644] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1208 ) );
  MX4XL \iRF_stage/reg_bank/U1204  ( .A(\iRF_stage/reg_bank/n1210 ), .B(
        \iRF_stage/reg_bank/n1208 ), .C(\iRF_stage/reg_bank/n1209 ), .D(
        \iRF_stage/reg_bank/n1207 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1211 ) );
  MX4X1 \iRF_stage/reg_bank/U1211  ( .A(\iRF_stage/reg_bank/reg_bank[613] ), 
        .B(\iRF_stage/reg_bank/reg_bank[581] ), .C(
        \iRF_stage/reg_bank/reg_bank[549] ), .D(
        \iRF_stage/reg_bank/reg_bank[517] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1217 ) );
  MX4X1 \iRF_stage/reg_bank/U1214  ( .A(\iRF_stage/reg_bank/reg_bank[997] ), 
        .B(\iRF_stage/reg_bank/reg_bank[965] ), .C(
        \iRF_stage/reg_bank/reg_bank[933] ), .D(
        \iRF_stage/reg_bank/reg_bank[901] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1220 ) );
  MX4X1 \iRF_stage/reg_bank/U1212  ( .A(\iRF_stage/reg_bank/reg_bank[741] ), 
        .B(\iRF_stage/reg_bank/reg_bank[709] ), .C(
        \iRF_stage/reg_bank/reg_bank[677] ), .D(
        \iRF_stage/reg_bank/reg_bank[645] ), .S0(n179), .S1(n204), .Y(
        \iRF_stage/reg_bank/n1218 ) );
  MX4XL \iRF_stage/reg_bank/U1215  ( .A(\iRF_stage/reg_bank/n1220 ), .B(
        \iRF_stage/reg_bank/n1218 ), .C(\iRF_stage/reg_bank/n1219 ), .D(
        \iRF_stage/reg_bank/n1217 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1221 ) );
  MX4X1 \iRF_stage/reg_bank/U1222  ( .A(\iRF_stage/reg_bank/reg_bank[614] ), 
        .B(\iRF_stage/reg_bank/reg_bank[582] ), .C(
        \iRF_stage/reg_bank/reg_bank[550] ), .D(
        \iRF_stage/reg_bank/reg_bank[518] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1227 ) );
  MX4X1 \iRF_stage/reg_bank/U1225  ( .A(\iRF_stage/reg_bank/reg_bank[998] ), 
        .B(\iRF_stage/reg_bank/reg_bank[966] ), .C(
        \iRF_stage/reg_bank/reg_bank[934] ), .D(
        \iRF_stage/reg_bank/reg_bank[902] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1230 ) );
  MX4X1 \iRF_stage/reg_bank/U1223  ( .A(\iRF_stage/reg_bank/reg_bank[742] ), 
        .B(\iRF_stage/reg_bank/reg_bank[710] ), .C(
        \iRF_stage/reg_bank/reg_bank[678] ), .D(
        \iRF_stage/reg_bank/reg_bank[646] ), .S0(n180), .S1(n205), .Y(
        \iRF_stage/reg_bank/n1228 ) );
  MX4XL \iRF_stage/reg_bank/U1226  ( .A(\iRF_stage/reg_bank/n1230 ), .B(
        \iRF_stage/reg_bank/n1228 ), .C(\iRF_stage/reg_bank/n1229 ), .D(
        \iRF_stage/reg_bank/n1227 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1231 ) );
  MX4X1 \iRF_stage/reg_bank/U1233  ( .A(\iRF_stage/reg_bank/reg_bank[615] ), 
        .B(\iRF_stage/reg_bank/reg_bank[583] ), .C(
        \iRF_stage/reg_bank/reg_bank[551] ), .D(
        \iRF_stage/reg_bank/reg_bank[519] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1237 ) );
  MX4X1 \iRF_stage/reg_bank/U1236  ( .A(\iRF_stage/reg_bank/reg_bank[999] ), 
        .B(\iRF_stage/reg_bank/reg_bank[967] ), .C(
        \iRF_stage/reg_bank/reg_bank[935] ), .D(
        \iRF_stage/reg_bank/reg_bank[903] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1240 ) );
  MX4X1 \iRF_stage/reg_bank/U1234  ( .A(\iRF_stage/reg_bank/reg_bank[743] ), 
        .B(\iRF_stage/reg_bank/reg_bank[711] ), .C(
        \iRF_stage/reg_bank/reg_bank[679] ), .D(
        \iRF_stage/reg_bank/reg_bank[647] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1238 ) );
  MX4XL \iRF_stage/reg_bank/U1237  ( .A(\iRF_stage/reg_bank/n1240 ), .B(
        \iRF_stage/reg_bank/n1238 ), .C(\iRF_stage/reg_bank/n1239 ), .D(
        \iRF_stage/reg_bank/n1237 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1241 ) );
  MX4X1 \iRF_stage/reg_bank/U1244  ( .A(\iRF_stage/reg_bank/reg_bank[616] ), 
        .B(\iRF_stage/reg_bank/reg_bank[584] ), .C(
        \iRF_stage/reg_bank/reg_bank[552] ), .D(
        \iRF_stage/reg_bank/reg_bank[520] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1247 ) );
  MX4X1 \iRF_stage/reg_bank/U1247  ( .A(\iRF_stage/reg_bank/reg_bank[1000] ), 
        .B(\iRF_stage/reg_bank/reg_bank[968] ), .C(
        \iRF_stage/reg_bank/reg_bank[936] ), .D(
        \iRF_stage/reg_bank/reg_bank[904] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1250 ) );
  MX4X1 \iRF_stage/reg_bank/U1245  ( .A(\iRF_stage/reg_bank/reg_bank[744] ), 
        .B(\iRF_stage/reg_bank/reg_bank[712] ), .C(
        \iRF_stage/reg_bank/reg_bank[680] ), .D(
        \iRF_stage/reg_bank/reg_bank[648] ), .S0(n181), .S1(n206), .Y(
        \iRF_stage/reg_bank/n1248 ) );
  MX4XL \iRF_stage/reg_bank/U1248  ( .A(\iRF_stage/reg_bank/n1250 ), .B(
        \iRF_stage/reg_bank/n1248 ), .C(\iRF_stage/reg_bank/n1249 ), .D(
        \iRF_stage/reg_bank/n1247 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1251 ) );
  MX4X1 \iRF_stage/reg_bank/U1255  ( .A(\iRF_stage/reg_bank/reg_bank[617] ), 
        .B(\iRF_stage/reg_bank/reg_bank[585] ), .C(
        \iRF_stage/reg_bank/reg_bank[553] ), .D(
        \iRF_stage/reg_bank/reg_bank[521] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1257 ) );
  MX4X1 \iRF_stage/reg_bank/U1258  ( .A(\iRF_stage/reg_bank/reg_bank[1001] ), 
        .B(\iRF_stage/reg_bank/reg_bank[969] ), .C(
        \iRF_stage/reg_bank/reg_bank[937] ), .D(
        \iRF_stage/reg_bank/reg_bank[905] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1260 ) );
  MX4X1 \iRF_stage/reg_bank/U1256  ( .A(\iRF_stage/reg_bank/reg_bank[745] ), 
        .B(\iRF_stage/reg_bank/reg_bank[713] ), .C(
        \iRF_stage/reg_bank/reg_bank[681] ), .D(
        \iRF_stage/reg_bank/reg_bank[649] ), .S0(n182), .S1(n207), .Y(
        \iRF_stage/reg_bank/n1258 ) );
  MX4XL \iRF_stage/reg_bank/U1259  ( .A(\iRF_stage/reg_bank/n1260 ), .B(
        \iRF_stage/reg_bank/n1258 ), .C(\iRF_stage/reg_bank/n1259 ), .D(
        \iRF_stage/reg_bank/n1257 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1261 ) );
  MX4X1 \iRF_stage/reg_bank/U1266  ( .A(\iRF_stage/reg_bank/reg_bank[618] ), 
        .B(\iRF_stage/reg_bank/reg_bank[586] ), .C(
        \iRF_stage/reg_bank/reg_bank[554] ), .D(
        \iRF_stage/reg_bank/reg_bank[522] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1267 ) );
  MX4X1 \iRF_stage/reg_bank/U1269  ( .A(\iRF_stage/reg_bank/reg_bank[1002] ), 
        .B(\iRF_stage/reg_bank/reg_bank[970] ), .C(
        \iRF_stage/reg_bank/reg_bank[938] ), .D(
        \iRF_stage/reg_bank/reg_bank[906] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1270 ) );
  MX4X1 \iRF_stage/reg_bank/U1267  ( .A(\iRF_stage/reg_bank/reg_bank[746] ), 
        .B(\iRF_stage/reg_bank/reg_bank[714] ), .C(
        \iRF_stage/reg_bank/reg_bank[682] ), .D(
        \iRF_stage/reg_bank/reg_bank[650] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1268 ) );
  MX4XL \iRF_stage/reg_bank/U1270  ( .A(\iRF_stage/reg_bank/n1270 ), .B(
        \iRF_stage/reg_bank/n1268 ), .C(\iRF_stage/reg_bank/n1269 ), .D(
        \iRF_stage/reg_bank/n1267 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1271 ) );
  MX4X1 \iRF_stage/reg_bank/U1277  ( .A(\iRF_stage/reg_bank/reg_bank[619] ), 
        .B(\iRF_stage/reg_bank/reg_bank[587] ), .C(
        \iRF_stage/reg_bank/reg_bank[555] ), .D(
        \iRF_stage/reg_bank/reg_bank[523] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1277 ) );
  MX4X1 \iRF_stage/reg_bank/U1280  ( .A(\iRF_stage/reg_bank/reg_bank[1003] ), 
        .B(\iRF_stage/reg_bank/reg_bank[971] ), .C(
        \iRF_stage/reg_bank/reg_bank[939] ), .D(
        \iRF_stage/reg_bank/reg_bank[907] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1280 ) );
  MX4X1 \iRF_stage/reg_bank/U1278  ( .A(\iRF_stage/reg_bank/reg_bank[747] ), 
        .B(\iRF_stage/reg_bank/reg_bank[715] ), .C(
        \iRF_stage/reg_bank/reg_bank[683] ), .D(
        \iRF_stage/reg_bank/reg_bank[651] ), .S0(n183), .S1(n208), .Y(
        \iRF_stage/reg_bank/n1278 ) );
  MX4XL \iRF_stage/reg_bank/U1281  ( .A(\iRF_stage/reg_bank/n1280 ), .B(
        \iRF_stage/reg_bank/n1278 ), .C(\iRF_stage/reg_bank/n1279 ), .D(
        \iRF_stage/reg_bank/n1277 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1281 ) );
  MX4X1 \iRF_stage/reg_bank/U1288  ( .A(\iRF_stage/reg_bank/reg_bank[620] ), 
        .B(\iRF_stage/reg_bank/reg_bank[588] ), .C(
        \iRF_stage/reg_bank/reg_bank[556] ), .D(
        \iRF_stage/reg_bank/reg_bank[524] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1287 ) );
  MX4X1 \iRF_stage/reg_bank/U1291  ( .A(\iRF_stage/reg_bank/reg_bank[1004] ), 
        .B(\iRF_stage/reg_bank/reg_bank[972] ), .C(
        \iRF_stage/reg_bank/reg_bank[940] ), .D(
        \iRF_stage/reg_bank/reg_bank[908] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1290 ) );
  MX4X1 \iRF_stage/reg_bank/U1289  ( .A(\iRF_stage/reg_bank/reg_bank[748] ), 
        .B(\iRF_stage/reg_bank/reg_bank[716] ), .C(
        \iRF_stage/reg_bank/reg_bank[684] ), .D(
        \iRF_stage/reg_bank/reg_bank[652] ), .S0(n184), .S1(n209), .Y(
        \iRF_stage/reg_bank/n1288 ) );
  MX4XL \iRF_stage/reg_bank/U1292  ( .A(\iRF_stage/reg_bank/n1290 ), .B(
        \iRF_stage/reg_bank/n1288 ), .C(\iRF_stage/reg_bank/n1289 ), .D(
        \iRF_stage/reg_bank/n1287 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1291 ) );
  MX4X1 \iRF_stage/reg_bank/U1299  ( .A(\iRF_stage/reg_bank/reg_bank[621] ), 
        .B(\iRF_stage/reg_bank/reg_bank[589] ), .C(
        \iRF_stage/reg_bank/reg_bank[557] ), .D(
        \iRF_stage/reg_bank/reg_bank[525] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1297 ) );
  MX4X1 \iRF_stage/reg_bank/U1302  ( .A(\iRF_stage/reg_bank/reg_bank[1005] ), 
        .B(\iRF_stage/reg_bank/reg_bank[973] ), .C(
        \iRF_stage/reg_bank/reg_bank[941] ), .D(
        \iRF_stage/reg_bank/reg_bank[909] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1300 ) );
  MX4X1 \iRF_stage/reg_bank/U1300  ( .A(\iRF_stage/reg_bank/reg_bank[749] ), 
        .B(\iRF_stage/reg_bank/reg_bank[717] ), .C(
        \iRF_stage/reg_bank/reg_bank[685] ), .D(
        \iRF_stage/reg_bank/reg_bank[653] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1298 ) );
  MX4XL \iRF_stage/reg_bank/U1303  ( .A(\iRF_stage/reg_bank/n1300 ), .B(
        \iRF_stage/reg_bank/n1298 ), .C(\iRF_stage/reg_bank/n1299 ), .D(
        \iRF_stage/reg_bank/n1297 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1301 ) );
  MX4X1 \iRF_stage/reg_bank/U1310  ( .A(\iRF_stage/reg_bank/reg_bank[622] ), 
        .B(\iRF_stage/reg_bank/reg_bank[590] ), .C(
        \iRF_stage/reg_bank/reg_bank[558] ), .D(
        \iRF_stage/reg_bank/reg_bank[526] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1307 ) );
  MX4X1 \iRF_stage/reg_bank/U1313  ( .A(\iRF_stage/reg_bank/reg_bank[1006] ), 
        .B(\iRF_stage/reg_bank/reg_bank[974] ), .C(
        \iRF_stage/reg_bank/reg_bank[942] ), .D(
        \iRF_stage/reg_bank/reg_bank[910] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1310 ) );
  MX4X1 \iRF_stage/reg_bank/U1311  ( .A(\iRF_stage/reg_bank/reg_bank[750] ), 
        .B(\iRF_stage/reg_bank/reg_bank[718] ), .C(
        \iRF_stage/reg_bank/reg_bank[686] ), .D(
        \iRF_stage/reg_bank/reg_bank[654] ), .S0(n185), .S1(n210), .Y(
        \iRF_stage/reg_bank/n1308 ) );
  MX4XL \iRF_stage/reg_bank/U1314  ( .A(\iRF_stage/reg_bank/n1310 ), .B(
        \iRF_stage/reg_bank/n1308 ), .C(\iRF_stage/reg_bank/n1309 ), .D(
        \iRF_stage/reg_bank/n1307 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1311 ) );
  MX4X1 \iRF_stage/reg_bank/U1321  ( .A(\iRF_stage/reg_bank/reg_bank[623] ), 
        .B(\iRF_stage/reg_bank/reg_bank[591] ), .C(
        \iRF_stage/reg_bank/reg_bank[559] ), .D(
        \iRF_stage/reg_bank/reg_bank[527] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1317 ) );
  MX4X1 \iRF_stage/reg_bank/U1324  ( .A(\iRF_stage/reg_bank/reg_bank[1007] ), 
        .B(\iRF_stage/reg_bank/reg_bank[975] ), .C(
        \iRF_stage/reg_bank/reg_bank[943] ), .D(
        \iRF_stage/reg_bank/reg_bank[911] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1320 ) );
  MX4X1 \iRF_stage/reg_bank/U1322  ( .A(\iRF_stage/reg_bank/reg_bank[751] ), 
        .B(\iRF_stage/reg_bank/reg_bank[719] ), .C(
        \iRF_stage/reg_bank/reg_bank[687] ), .D(
        \iRF_stage/reg_bank/reg_bank[655] ), .S0(n186), .S1(n211), .Y(
        \iRF_stage/reg_bank/n1318 ) );
  MX4XL \iRF_stage/reg_bank/U1325  ( .A(\iRF_stage/reg_bank/n1320 ), .B(
        \iRF_stage/reg_bank/n1318 ), .C(\iRF_stage/reg_bank/n1319 ), .D(
        \iRF_stage/reg_bank/n1317 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1321 ) );
  MX4X1 \iRF_stage/reg_bank/U1332  ( .A(\iRF_stage/reg_bank/reg_bank[624] ), 
        .B(\iRF_stage/reg_bank/reg_bank[592] ), .C(
        \iRF_stage/reg_bank/reg_bank[560] ), .D(
        \iRF_stage/reg_bank/reg_bank[528] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1327 ) );
  MX4X1 \iRF_stage/reg_bank/U1335  ( .A(\iRF_stage/reg_bank/reg_bank[1008] ), 
        .B(\iRF_stage/reg_bank/reg_bank[976] ), .C(
        \iRF_stage/reg_bank/reg_bank[944] ), .D(
        \iRF_stage/reg_bank/reg_bank[912] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1330 ) );
  MX4X1 \iRF_stage/reg_bank/U1333  ( .A(\iRF_stage/reg_bank/reg_bank[752] ), 
        .B(\iRF_stage/reg_bank/reg_bank[720] ), .C(
        \iRF_stage/reg_bank/reg_bank[688] ), .D(
        \iRF_stage/reg_bank/reg_bank[656] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1328 ) );
  MX4XL \iRF_stage/reg_bank/U1336  ( .A(\iRF_stage/reg_bank/n1330 ), .B(
        \iRF_stage/reg_bank/n1328 ), .C(\iRF_stage/reg_bank/n1329 ), .D(
        \iRF_stage/reg_bank/n1327 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1331 ) );
  MX4X1 \iRF_stage/reg_bank/U1343  ( .A(\iRF_stage/reg_bank/reg_bank[625] ), 
        .B(\iRF_stage/reg_bank/reg_bank[593] ), .C(
        \iRF_stage/reg_bank/reg_bank[561] ), .D(
        \iRF_stage/reg_bank/reg_bank[529] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1337 ) );
  MX4X1 \iRF_stage/reg_bank/U1346  ( .A(\iRF_stage/reg_bank/reg_bank[1009] ), 
        .B(\iRF_stage/reg_bank/reg_bank[977] ), .C(
        \iRF_stage/reg_bank/reg_bank[945] ), .D(
        \iRF_stage/reg_bank/reg_bank[913] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1340 ) );
  MX4X1 \iRF_stage/reg_bank/U1344  ( .A(\iRF_stage/reg_bank/reg_bank[753] ), 
        .B(\iRF_stage/reg_bank/reg_bank[721] ), .C(
        \iRF_stage/reg_bank/reg_bank[689] ), .D(
        \iRF_stage/reg_bank/reg_bank[657] ), .S0(n187), .S1(n212), .Y(
        \iRF_stage/reg_bank/n1338 ) );
  MX4XL \iRF_stage/reg_bank/U1347  ( .A(\iRF_stage/reg_bank/n1340 ), .B(
        \iRF_stage/reg_bank/n1338 ), .C(\iRF_stage/reg_bank/n1339 ), .D(
        \iRF_stage/reg_bank/n1337 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1341 ) );
  MX4X1 \iRF_stage/reg_bank/U1354  ( .A(\iRF_stage/reg_bank/reg_bank[626] ), 
        .B(\iRF_stage/reg_bank/reg_bank[594] ), .C(
        \iRF_stage/reg_bank/reg_bank[562] ), .D(
        \iRF_stage/reg_bank/reg_bank[530] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1347 ) );
  MX4X1 \iRF_stage/reg_bank/U1357  ( .A(\iRF_stage/reg_bank/reg_bank[1010] ), 
        .B(\iRF_stage/reg_bank/reg_bank[978] ), .C(
        \iRF_stage/reg_bank/reg_bank[946] ), .D(
        \iRF_stage/reg_bank/reg_bank[914] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1350 ) );
  MX4X1 \iRF_stage/reg_bank/U1355  ( .A(\iRF_stage/reg_bank/reg_bank[754] ), 
        .B(\iRF_stage/reg_bank/reg_bank[722] ), .C(
        \iRF_stage/reg_bank/reg_bank[690] ), .D(
        \iRF_stage/reg_bank/reg_bank[658] ), .S0(n188), .S1(n213), .Y(
        \iRF_stage/reg_bank/n1348 ) );
  MX4XL \iRF_stage/reg_bank/U1358  ( .A(\iRF_stage/reg_bank/n1350 ), .B(
        \iRF_stage/reg_bank/n1348 ), .C(\iRF_stage/reg_bank/n1349 ), .D(
        \iRF_stage/reg_bank/n1347 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1351 ) );
  MX4X1 \iRF_stage/reg_bank/U1365  ( .A(\iRF_stage/reg_bank/reg_bank[627] ), 
        .B(\iRF_stage/reg_bank/reg_bank[595] ), .C(
        \iRF_stage/reg_bank/reg_bank[563] ), .D(
        \iRF_stage/reg_bank/reg_bank[531] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1357 ) );
  MX4X1 \iRF_stage/reg_bank/U1368  ( .A(\iRF_stage/reg_bank/reg_bank[1011] ), 
        .B(\iRF_stage/reg_bank/reg_bank[979] ), .C(
        \iRF_stage/reg_bank/reg_bank[947] ), .D(
        \iRF_stage/reg_bank/reg_bank[915] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1360 ) );
  MX4X1 \iRF_stage/reg_bank/U1366  ( .A(\iRF_stage/reg_bank/reg_bank[755] ), 
        .B(\iRF_stage/reg_bank/reg_bank[723] ), .C(
        \iRF_stage/reg_bank/reg_bank[691] ), .D(
        \iRF_stage/reg_bank/reg_bank[659] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1358 ) );
  MX4XL \iRF_stage/reg_bank/U1369  ( .A(\iRF_stage/reg_bank/n1360 ), .B(
        \iRF_stage/reg_bank/n1358 ), .C(\iRF_stage/reg_bank/n1359 ), .D(
        \iRF_stage/reg_bank/n1357 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1361 ) );
  MX4X1 \iRF_stage/reg_bank/U1376  ( .A(\iRF_stage/reg_bank/reg_bank[628] ), 
        .B(\iRF_stage/reg_bank/reg_bank[596] ), .C(
        \iRF_stage/reg_bank/reg_bank[564] ), .D(
        \iRF_stage/reg_bank/reg_bank[532] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1367 ) );
  MX4X1 \iRF_stage/reg_bank/U1379  ( .A(\iRF_stage/reg_bank/reg_bank[1012] ), 
        .B(\iRF_stage/reg_bank/reg_bank[980] ), .C(
        \iRF_stage/reg_bank/reg_bank[948] ), .D(
        \iRF_stage/reg_bank/reg_bank[916] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1370 ) );
  MX4X1 \iRF_stage/reg_bank/U1377  ( .A(\iRF_stage/reg_bank/reg_bank[756] ), 
        .B(\iRF_stage/reg_bank/reg_bank[724] ), .C(
        \iRF_stage/reg_bank/reg_bank[692] ), .D(
        \iRF_stage/reg_bank/reg_bank[660] ), .S0(n189), .S1(n214), .Y(
        \iRF_stage/reg_bank/n1368 ) );
  MX4XL \iRF_stage/reg_bank/U1380  ( .A(\iRF_stage/reg_bank/n1370 ), .B(
        \iRF_stage/reg_bank/n1368 ), .C(\iRF_stage/reg_bank/n1369 ), .D(
        \iRF_stage/reg_bank/n1367 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1371 ) );
  MX4X1 \iRF_stage/reg_bank/U1387  ( .A(\iRF_stage/reg_bank/reg_bank[629] ), 
        .B(\iRF_stage/reg_bank/reg_bank[597] ), .C(
        \iRF_stage/reg_bank/reg_bank[565] ), .D(
        \iRF_stage/reg_bank/reg_bank[533] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1377 ) );
  MX4X1 \iRF_stage/reg_bank/U1390  ( .A(\iRF_stage/reg_bank/reg_bank[1013] ), 
        .B(\iRF_stage/reg_bank/reg_bank[981] ), .C(
        \iRF_stage/reg_bank/reg_bank[949] ), .D(
        \iRF_stage/reg_bank/reg_bank[917] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1380 ) );
  MX4X1 \iRF_stage/reg_bank/U1388  ( .A(\iRF_stage/reg_bank/reg_bank[757] ), 
        .B(\iRF_stage/reg_bank/reg_bank[725] ), .C(
        \iRF_stage/reg_bank/reg_bank[693] ), .D(
        \iRF_stage/reg_bank/reg_bank[661] ), .S0(n190), .S1(n215), .Y(
        \iRF_stage/reg_bank/n1378 ) );
  MX4XL \iRF_stage/reg_bank/U1391  ( .A(\iRF_stage/reg_bank/n1380 ), .B(
        \iRF_stage/reg_bank/n1378 ), .C(\iRF_stage/reg_bank/n1379 ), .D(
        \iRF_stage/reg_bank/n1377 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1381 ) );
  MX4X1 \iRF_stage/reg_bank/U1398  ( .A(\iRF_stage/reg_bank/reg_bank[630] ), 
        .B(\iRF_stage/reg_bank/reg_bank[598] ), .C(
        \iRF_stage/reg_bank/reg_bank[566] ), .D(
        \iRF_stage/reg_bank/reg_bank[534] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1387 ) );
  MX4X1 \iRF_stage/reg_bank/U1401  ( .A(\iRF_stage/reg_bank/reg_bank[1014] ), 
        .B(\iRF_stage/reg_bank/reg_bank[982] ), .C(
        \iRF_stage/reg_bank/reg_bank[950] ), .D(
        \iRF_stage/reg_bank/reg_bank[918] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1390 ) );
  MX4X1 \iRF_stage/reg_bank/U1399  ( .A(\iRF_stage/reg_bank/reg_bank[758] ), 
        .B(\iRF_stage/reg_bank/reg_bank[726] ), .C(
        \iRF_stage/reg_bank/reg_bank[694] ), .D(
        \iRF_stage/reg_bank/reg_bank[662] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1388 ) );
  MX4XL \iRF_stage/reg_bank/U1402  ( .A(\iRF_stage/reg_bank/n1390 ), .B(
        \iRF_stage/reg_bank/n1388 ), .C(\iRF_stage/reg_bank/n1389 ), .D(
        \iRF_stage/reg_bank/n1387 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1391 ) );
  MX4X1 \iRF_stage/reg_bank/U1409  ( .A(\iRF_stage/reg_bank/reg_bank[631] ), 
        .B(\iRF_stage/reg_bank/reg_bank[599] ), .C(
        \iRF_stage/reg_bank/reg_bank[567] ), .D(
        \iRF_stage/reg_bank/reg_bank[535] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1397 ) );
  MX4X1 \iRF_stage/reg_bank/U1412  ( .A(\iRF_stage/reg_bank/reg_bank[1015] ), 
        .B(\iRF_stage/reg_bank/reg_bank[983] ), .C(
        \iRF_stage/reg_bank/reg_bank[951] ), .D(
        \iRF_stage/reg_bank/reg_bank[919] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1400 ) );
  MX4X1 \iRF_stage/reg_bank/U1410  ( .A(\iRF_stage/reg_bank/reg_bank[759] ), 
        .B(\iRF_stage/reg_bank/reg_bank[727] ), .C(
        \iRF_stage/reg_bank/reg_bank[695] ), .D(
        \iRF_stage/reg_bank/reg_bank[663] ), .S0(n191), .S1(n216), .Y(
        \iRF_stage/reg_bank/n1398 ) );
  MX4XL \iRF_stage/reg_bank/U1413  ( .A(\iRF_stage/reg_bank/n1400 ), .B(
        \iRF_stage/reg_bank/n1398 ), .C(\iRF_stage/reg_bank/n1399 ), .D(
        \iRF_stage/reg_bank/n1397 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1401 ) );
  MX4X1 \iRF_stage/reg_bank/U1420  ( .A(\iRF_stage/reg_bank/reg_bank[632] ), 
        .B(\iRF_stage/reg_bank/reg_bank[600] ), .C(
        \iRF_stage/reg_bank/reg_bank[568] ), .D(
        \iRF_stage/reg_bank/reg_bank[536] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1407 ) );
  MX4X1 \iRF_stage/reg_bank/U1423  ( .A(\iRF_stage/reg_bank/reg_bank[1016] ), 
        .B(\iRF_stage/reg_bank/reg_bank[984] ), .C(
        \iRF_stage/reg_bank/reg_bank[952] ), .D(
        \iRF_stage/reg_bank/reg_bank[920] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1410 ) );
  MX4X1 \iRF_stage/reg_bank/U1421  ( .A(\iRF_stage/reg_bank/reg_bank[760] ), 
        .B(\iRF_stage/reg_bank/reg_bank[728] ), .C(
        \iRF_stage/reg_bank/reg_bank[696] ), .D(
        \iRF_stage/reg_bank/reg_bank[664] ), .S0(n192), .S1(n217), .Y(
        \iRF_stage/reg_bank/n1408 ) );
  MX4XL \iRF_stage/reg_bank/U1424  ( .A(\iRF_stage/reg_bank/n1410 ), .B(
        \iRF_stage/reg_bank/n1408 ), .C(\iRF_stage/reg_bank/n1409 ), .D(
        \iRF_stage/reg_bank/n1407 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1411 ) );
  MX4X1 \iRF_stage/reg_bank/U1431  ( .A(\iRF_stage/reg_bank/reg_bank[633] ), 
        .B(\iRF_stage/reg_bank/reg_bank[601] ), .C(
        \iRF_stage/reg_bank/reg_bank[569] ), .D(
        \iRF_stage/reg_bank/reg_bank[537] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1417 ) );
  MX4X1 \iRF_stage/reg_bank/U1434  ( .A(\iRF_stage/reg_bank/reg_bank[1017] ), 
        .B(\iRF_stage/reg_bank/reg_bank[985] ), .C(
        \iRF_stage/reg_bank/reg_bank[953] ), .D(
        \iRF_stage/reg_bank/reg_bank[921] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1420 ) );
  MX4X1 \iRF_stage/reg_bank/U1432  ( .A(\iRF_stage/reg_bank/reg_bank[761] ), 
        .B(\iRF_stage/reg_bank/reg_bank[729] ), .C(
        \iRF_stage/reg_bank/reg_bank[697] ), .D(
        \iRF_stage/reg_bank/reg_bank[665] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1418 ) );
  MX4XL \iRF_stage/reg_bank/U1435  ( .A(\iRF_stage/reg_bank/n1420 ), .B(
        \iRF_stage/reg_bank/n1418 ), .C(\iRF_stage/reg_bank/n1419 ), .D(
        \iRF_stage/reg_bank/n1417 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1421 ) );
  MX4X1 \iRF_stage/reg_bank/U1442  ( .A(\iRF_stage/reg_bank/reg_bank[634] ), 
        .B(\iRF_stage/reg_bank/reg_bank[602] ), .C(
        \iRF_stage/reg_bank/reg_bank[570] ), .D(
        \iRF_stage/reg_bank/reg_bank[538] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1427 ) );
  MX4X1 \iRF_stage/reg_bank/U1445  ( .A(\iRF_stage/reg_bank/reg_bank[1018] ), 
        .B(\iRF_stage/reg_bank/reg_bank[986] ), .C(
        \iRF_stage/reg_bank/reg_bank[954] ), .D(
        \iRF_stage/reg_bank/reg_bank[922] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1430 ) );
  MX4X1 \iRF_stage/reg_bank/U1443  ( .A(\iRF_stage/reg_bank/reg_bank[762] ), 
        .B(\iRF_stage/reg_bank/reg_bank[730] ), .C(
        \iRF_stage/reg_bank/reg_bank[698] ), .D(
        \iRF_stage/reg_bank/reg_bank[666] ), .S0(n193), .S1(n218), .Y(
        \iRF_stage/reg_bank/n1428 ) );
  MX4XL \iRF_stage/reg_bank/U1446  ( .A(\iRF_stage/reg_bank/n1430 ), .B(
        \iRF_stage/reg_bank/n1428 ), .C(\iRF_stage/reg_bank/n1429 ), .D(
        \iRF_stage/reg_bank/n1427 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1431 ) );
  MX4X1 \iRF_stage/reg_bank/U1453  ( .A(\iRF_stage/reg_bank/reg_bank[635] ), 
        .B(\iRF_stage/reg_bank/reg_bank[603] ), .C(
        \iRF_stage/reg_bank/reg_bank[571] ), .D(
        \iRF_stage/reg_bank/reg_bank[539] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1437 ) );
  MX4X1 \iRF_stage/reg_bank/U1456  ( .A(\iRF_stage/reg_bank/reg_bank[1019] ), 
        .B(\iRF_stage/reg_bank/reg_bank[987] ), .C(
        \iRF_stage/reg_bank/reg_bank[955] ), .D(
        \iRF_stage/reg_bank/reg_bank[923] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1440 ) );
  MX4X1 \iRF_stage/reg_bank/U1454  ( .A(\iRF_stage/reg_bank/reg_bank[763] ), 
        .B(\iRF_stage/reg_bank/reg_bank[731] ), .C(
        \iRF_stage/reg_bank/reg_bank[699] ), .D(
        \iRF_stage/reg_bank/reg_bank[667] ), .S0(n194), .S1(n219), .Y(
        \iRF_stage/reg_bank/n1438 ) );
  MX4XL \iRF_stage/reg_bank/U1457  ( .A(\iRF_stage/reg_bank/n1440 ), .B(
        \iRF_stage/reg_bank/n1438 ), .C(\iRF_stage/reg_bank/n1439 ), .D(
        \iRF_stage/reg_bank/n1437 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1441 ) );
  MX4X1 \iRF_stage/reg_bank/U1464  ( .A(\iRF_stage/reg_bank/reg_bank[636] ), 
        .B(\iRF_stage/reg_bank/reg_bank[604] ), .C(
        \iRF_stage/reg_bank/reg_bank[572] ), .D(
        \iRF_stage/reg_bank/reg_bank[540] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1447 ) );
  MX4X1 \iRF_stage/reg_bank/U1467  ( .A(\iRF_stage/reg_bank/reg_bank[1020] ), 
        .B(\iRF_stage/reg_bank/reg_bank[988] ), .C(
        \iRF_stage/reg_bank/reg_bank[956] ), .D(
        \iRF_stage/reg_bank/reg_bank[924] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1450 ) );
  MX4X1 \iRF_stage/reg_bank/U1465  ( .A(\iRF_stage/reg_bank/reg_bank[764] ), 
        .B(\iRF_stage/reg_bank/reg_bank[732] ), .C(
        \iRF_stage/reg_bank/reg_bank[700] ), .D(
        \iRF_stage/reg_bank/reg_bank[668] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1448 ) );
  MX4XL \iRF_stage/reg_bank/U1468  ( .A(\iRF_stage/reg_bank/n1450 ), .B(
        \iRF_stage/reg_bank/n1448 ), .C(\iRF_stage/reg_bank/n1449 ), .D(
        \iRF_stage/reg_bank/n1447 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1451 ) );
  MX4X1 \iRF_stage/reg_bank/U1475  ( .A(\iRF_stage/reg_bank/reg_bank[637] ), 
        .B(\iRF_stage/reg_bank/reg_bank[605] ), .C(
        \iRF_stage/reg_bank/reg_bank[573] ), .D(
        \iRF_stage/reg_bank/reg_bank[541] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1457 ) );
  MX4X1 \iRF_stage/reg_bank/U1478  ( .A(\iRF_stage/reg_bank/reg_bank[1021] ), 
        .B(\iRF_stage/reg_bank/reg_bank[989] ), .C(
        \iRF_stage/reg_bank/reg_bank[957] ), .D(
        \iRF_stage/reg_bank/reg_bank[925] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1460 ) );
  MX4X1 \iRF_stage/reg_bank/U1476  ( .A(\iRF_stage/reg_bank/reg_bank[765] ), 
        .B(\iRF_stage/reg_bank/reg_bank[733] ), .C(
        \iRF_stage/reg_bank/reg_bank[701] ), .D(
        \iRF_stage/reg_bank/reg_bank[669] ), .S0(n195), .S1(n220), .Y(
        \iRF_stage/reg_bank/n1458 ) );
  MX4XL \iRF_stage/reg_bank/U1479  ( .A(\iRF_stage/reg_bank/n1460 ), .B(
        \iRF_stage/reg_bank/n1458 ), .C(\iRF_stage/reg_bank/n1459 ), .D(
        \iRF_stage/reg_bank/n1457 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1461 ) );
  MX4X1 \iRF_stage/reg_bank/U1486  ( .A(\iRF_stage/reg_bank/reg_bank[638] ), 
        .B(\iRF_stage/reg_bank/reg_bank[606] ), .C(
        \iRF_stage/reg_bank/reg_bank[574] ), .D(
        \iRF_stage/reg_bank/reg_bank[542] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1467 ) );
  MX4X1 \iRF_stage/reg_bank/U1489  ( .A(\iRF_stage/reg_bank/reg_bank[1022] ), 
        .B(\iRF_stage/reg_bank/reg_bank[990] ), .C(
        \iRF_stage/reg_bank/reg_bank[958] ), .D(
        \iRF_stage/reg_bank/reg_bank[926] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1470 ) );
  MX4X1 \iRF_stage/reg_bank/U1487  ( .A(\iRF_stage/reg_bank/reg_bank[766] ), 
        .B(\iRF_stage/reg_bank/reg_bank[734] ), .C(
        \iRF_stage/reg_bank/reg_bank[702] ), .D(
        \iRF_stage/reg_bank/reg_bank[670] ), .S0(n196), .S1(n221), .Y(
        \iRF_stage/reg_bank/n1468 ) );
  MX4XL \iRF_stage/reg_bank/U1490  ( .A(\iRF_stage/reg_bank/n1470 ), .B(
        \iRF_stage/reg_bank/n1468 ), .C(\iRF_stage/reg_bank/n1469 ), .D(
        \iRF_stage/reg_bank/n1467 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1471 ) );
  MX4X1 \iRF_stage/reg_bank/U1497  ( .A(\iRF_stage/reg_bank/reg_bank[639] ), 
        .B(\iRF_stage/reg_bank/reg_bank[607] ), .C(
        \iRF_stage/reg_bank/reg_bank[575] ), .D(
        \iRF_stage/reg_bank/reg_bank[543] ), .S0(n197), .S1(
        \iRF_stage/reg_bank/N13 ), .Y(\iRF_stage/reg_bank/n1477 ) );
  MX4X1 \iRF_stage/reg_bank/U1500  ( .A(\iRF_stage/reg_bank/reg_bank[1023] ), 
        .B(\iRF_stage/reg_bank/reg_bank[991] ), .C(
        \iRF_stage/reg_bank/reg_bank[959] ), .D(
        \iRF_stage/reg_bank/reg_bank[927] ), .S0(n197), .S1(
        \iRF_stage/reg_bank/N13 ), .Y(\iRF_stage/reg_bank/n1480 ) );
  MX4X1 \iRF_stage/reg_bank/U1498  ( .A(\iRF_stage/reg_bank/reg_bank[767] ), 
        .B(\iRF_stage/reg_bank/reg_bank[735] ), .C(
        \iRF_stage/reg_bank/reg_bank[703] ), .D(
        \iRF_stage/reg_bank/reg_bank[671] ), .S0(n197), .S1(
        \iRF_stage/reg_bank/N13 ), .Y(\iRF_stage/reg_bank/n1478 ) );
  MX4X1 \iRF_stage/reg_bank/U1501  ( .A(\iRF_stage/reg_bank/n1480 ), .B(
        \iRF_stage/reg_bank/n1478 ), .C(\iRF_stage/reg_bank/n1479 ), .D(
        \iRF_stage/reg_bank/n1477 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1481 ) );
  XOR3X2 \iRF_stage/i_pc_gen/r62/U1_31  ( .A(BUS27031[31]), .B(1'b0), .C(
        \iRF_stage/i_pc_gen/r62/carry[31] ), .Y(\iRF_stage/i_pc_gen/N65 ) );
  MX4XL \iRF_stage/reg_bank/U1507  ( .A(\iRF_stage/reg_bank/n1485 ), .B(
        \iRF_stage/reg_bank/n1483 ), .C(\iRF_stage/reg_bank/n1484 ), .D(
        \iRF_stage/reg_bank/n1482 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1486 ) );
  MX2X2 \iRF_stage/reg_bank/U1513  ( .A(\iRF_stage/reg_bank/n1491 ), .B(
        \iRF_stage/reg_bank/n1486 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1120 ) );
  MX4XL \iRF_stage/reg_bank/U1529  ( .A(\iRF_stage/reg_bank/n1505 ), .B(
        \iRF_stage/reg_bank/n1503 ), .C(\iRF_stage/reg_bank/n1504 ), .D(
        \iRF_stage/reg_bank/n1502 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1506 ) );
  MX2X2 \iRF_stage/reg_bank/U1535  ( .A(\iRF_stage/reg_bank/n1511 ), .B(
        \iRF_stage/reg_bank/n1506 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1118 ) );
  MX4X1 \iRF_stage/reg_bank/U1617  ( .A(\iRF_stage/reg_bank/n1585 ), .B(
        \iRF_stage/reg_bank/n1583 ), .C(\iRF_stage/reg_bank/n1584 ), .D(
        \iRF_stage/reg_bank/n1582 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1586 ) );
  MX2X2 \iRF_stage/reg_bank/U1623  ( .A(\iRF_stage/reg_bank/n1591 ), .B(
        \iRF_stage/reg_bank/n1586 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1110 ) );
  MX4X1 \iRF_stage/reg_bank/U1628  ( .A(\iRF_stage/reg_bank/n1595 ), .B(
        \iRF_stage/reg_bank/n1593 ), .C(\iRF_stage/reg_bank/n1594 ), .D(
        \iRF_stage/reg_bank/n1592 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1596 ) );
  MX2X2 \iRF_stage/reg_bank/U1634  ( .A(\iRF_stage/reg_bank/n1601 ), .B(
        \iRF_stage/reg_bank/n1596 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1109 ) );
  MX4X1 \iRF_stage/reg_bank/U1848  ( .A(\iRF_stage/reg_bank/n1795 ), .B(
        \iRF_stage/reg_bank/n1793 ), .C(\iRF_stage/reg_bank/n1794 ), .D(
        \iRF_stage/reg_bank/n1792 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1796 ) );
  MX2X2 \iRF_stage/reg_bank/U1854  ( .A(\iRF_stage/reg_bank/n1801 ), .B(
        \iRF_stage/reg_bank/n1796 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1089 ) );
  MX4X1 \iRF_stage/reg_bank/U1518  ( .A(\iRF_stage/reg_bank/n1495 ), .B(
        \iRF_stage/reg_bank/n1493 ), .C(\iRF_stage/reg_bank/n1494 ), .D(
        \iRF_stage/reg_bank/n1492 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1496 ) );
  MX2X2 \iRF_stage/reg_bank/U1524  ( .A(\iRF_stage/reg_bank/n1501 ), .B(
        \iRF_stage/reg_bank/n1496 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1119 ) );
  MX4X1 \iRF_stage/reg_bank/U1540  ( .A(\iRF_stage/reg_bank/n1515 ), .B(
        \iRF_stage/reg_bank/n1513 ), .C(\iRF_stage/reg_bank/n1514 ), .D(
        \iRF_stage/reg_bank/n1512 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1516 ) );
  MX2X2 \iRF_stage/reg_bank/U1546  ( .A(\iRF_stage/reg_bank/n1521 ), .B(
        \iRF_stage/reg_bank/n1516 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1117 ) );
  MX4X1 \iRF_stage/reg_bank/U1551  ( .A(\iRF_stage/reg_bank/n1525 ), .B(
        \iRF_stage/reg_bank/n1523 ), .C(\iRF_stage/reg_bank/n1524 ), .D(
        \iRF_stage/reg_bank/n1522 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1526 ) );
  MX2X2 \iRF_stage/reg_bank/U1557  ( .A(\iRF_stage/reg_bank/n1531 ), .B(
        \iRF_stage/reg_bank/n1526 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1116 ) );
  MX4X1 \iRF_stage/reg_bank/U1562  ( .A(\iRF_stage/reg_bank/n1535 ), .B(
        \iRF_stage/reg_bank/n1533 ), .C(\iRF_stage/reg_bank/n1534 ), .D(
        \iRF_stage/reg_bank/n1532 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1536 ) );
  MX2X2 \iRF_stage/reg_bank/U1568  ( .A(\iRF_stage/reg_bank/n1541 ), .B(
        \iRF_stage/reg_bank/n1536 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1115 ) );
  MX4X1 \iRF_stage/reg_bank/U1573  ( .A(\iRF_stage/reg_bank/n1545 ), .B(
        \iRF_stage/reg_bank/n1543 ), .C(\iRF_stage/reg_bank/n1544 ), .D(
        \iRF_stage/reg_bank/n1542 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1546 ) );
  MX2X2 \iRF_stage/reg_bank/U1579  ( .A(\iRF_stage/reg_bank/n1551 ), .B(
        \iRF_stage/reg_bank/n1546 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1114 ) );
  MX4X1 \iRF_stage/reg_bank/U1584  ( .A(\iRF_stage/reg_bank/n1555 ), .B(
        \iRF_stage/reg_bank/n1553 ), .C(\iRF_stage/reg_bank/n1554 ), .D(
        \iRF_stage/reg_bank/n1552 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1556 ) );
  MX2X2 \iRF_stage/reg_bank/U1590  ( .A(\iRF_stage/reg_bank/n1561 ), .B(
        \iRF_stage/reg_bank/n1556 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1113 ) );
  MX4X1 \iRF_stage/reg_bank/U1595  ( .A(\iRF_stage/reg_bank/n1565 ), .B(
        \iRF_stage/reg_bank/n1563 ), .C(\iRF_stage/reg_bank/n1564 ), .D(
        \iRF_stage/reg_bank/n1562 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1566 ) );
  MX2X2 \iRF_stage/reg_bank/U1601  ( .A(\iRF_stage/reg_bank/n1571 ), .B(
        \iRF_stage/reg_bank/n1566 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1112 ) );
  MX4X1 \iRF_stage/reg_bank/U1606  ( .A(\iRF_stage/reg_bank/n1575 ), .B(
        \iRF_stage/reg_bank/n1573 ), .C(\iRF_stage/reg_bank/n1574 ), .D(
        \iRF_stage/reg_bank/n1572 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1576 ) );
  MX2X2 \iRF_stage/reg_bank/U1612  ( .A(\iRF_stage/reg_bank/n1581 ), .B(
        \iRF_stage/reg_bank/n1576 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1111 ) );
  MX4X1 \iRF_stage/reg_bank/U1639  ( .A(\iRF_stage/reg_bank/n1605 ), .B(
        \iRF_stage/reg_bank/n1603 ), .C(\iRF_stage/reg_bank/n1604 ), .D(
        \iRF_stage/reg_bank/n1602 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1606 ) );
  MX2X2 \iRF_stage/reg_bank/U1645  ( .A(\iRF_stage/reg_bank/n1611 ), .B(
        \iRF_stage/reg_bank/n1606 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1108 ) );
  MX4X1 \iRF_stage/reg_bank/U1650  ( .A(\iRF_stage/reg_bank/n1615 ), .B(
        \iRF_stage/reg_bank/n1613 ), .C(\iRF_stage/reg_bank/n1614 ), .D(
        \iRF_stage/reg_bank/n1612 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1616 ) );
  MX2X2 \iRF_stage/reg_bank/U1656  ( .A(\iRF_stage/reg_bank/n1621 ), .B(
        \iRF_stage/reg_bank/n1616 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1107 ) );
  MX4X1 \iRF_stage/reg_bank/U1661  ( .A(\iRF_stage/reg_bank/n1625 ), .B(
        \iRF_stage/reg_bank/n1623 ), .C(\iRF_stage/reg_bank/n1624 ), .D(
        \iRF_stage/reg_bank/n1622 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1626 ) );
  MX2X2 \iRF_stage/reg_bank/U1667  ( .A(\iRF_stage/reg_bank/n1631 ), .B(
        \iRF_stage/reg_bank/n1626 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1106 ) );
  MX4X1 \iRF_stage/reg_bank/U1672  ( .A(\iRF_stage/reg_bank/n1635 ), .B(
        \iRF_stage/reg_bank/n1633 ), .C(\iRF_stage/reg_bank/n1634 ), .D(
        \iRF_stage/reg_bank/n1632 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1636 ) );
  MX2X2 \iRF_stage/reg_bank/U1678  ( .A(\iRF_stage/reg_bank/n1641 ), .B(
        \iRF_stage/reg_bank/n1636 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1105 ) );
  MX4X1 \iRF_stage/reg_bank/U1683  ( .A(\iRF_stage/reg_bank/n1645 ), .B(
        \iRF_stage/reg_bank/n1643 ), .C(\iRF_stage/reg_bank/n1644 ), .D(
        \iRF_stage/reg_bank/n1642 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1646 ) );
  MX2X2 \iRF_stage/reg_bank/U1689  ( .A(\iRF_stage/reg_bank/n1651 ), .B(
        \iRF_stage/reg_bank/n1646 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1104 ) );
  MX4X1 \iRF_stage/reg_bank/U1694  ( .A(\iRF_stage/reg_bank/n1655 ), .B(
        \iRF_stage/reg_bank/n1653 ), .C(\iRF_stage/reg_bank/n1654 ), .D(
        \iRF_stage/reg_bank/n1652 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1656 ) );
  MX2X2 \iRF_stage/reg_bank/U1700  ( .A(\iRF_stage/reg_bank/n1661 ), .B(
        \iRF_stage/reg_bank/n1656 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1103 ) );
  MX4X1 \iRF_stage/reg_bank/U1705  ( .A(\iRF_stage/reg_bank/n1665 ), .B(
        \iRF_stage/reg_bank/n1663 ), .C(\iRF_stage/reg_bank/n1664 ), .D(
        \iRF_stage/reg_bank/n1662 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1666 ) );
  MX2X2 \iRF_stage/reg_bank/U1711  ( .A(\iRF_stage/reg_bank/n1671 ), .B(
        \iRF_stage/reg_bank/n1666 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1102 ) );
  MX4X1 \iRF_stage/reg_bank/U1716  ( .A(\iRF_stage/reg_bank/n1675 ), .B(
        \iRF_stage/reg_bank/n1673 ), .C(\iRF_stage/reg_bank/n1674 ), .D(
        \iRF_stage/reg_bank/n1672 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1676 ) );
  MX2X2 \iRF_stage/reg_bank/U1722  ( .A(\iRF_stage/reg_bank/n1681 ), .B(
        \iRF_stage/reg_bank/n1676 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1101 ) );
  MX4X1 \iRF_stage/reg_bank/U1727  ( .A(\iRF_stage/reg_bank/n1685 ), .B(
        \iRF_stage/reg_bank/n1683 ), .C(\iRF_stage/reg_bank/n1684 ), .D(
        \iRF_stage/reg_bank/n1682 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1686 ) );
  MX2X2 \iRF_stage/reg_bank/U1733  ( .A(\iRF_stage/reg_bank/n1691 ), .B(
        \iRF_stage/reg_bank/n1686 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1100 ) );
  MX4X1 \iRF_stage/reg_bank/U1738  ( .A(\iRF_stage/reg_bank/n1695 ), .B(
        \iRF_stage/reg_bank/n1693 ), .C(\iRF_stage/reg_bank/n1694 ), .D(
        \iRF_stage/reg_bank/n1692 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1696 ) );
  MX2X2 \iRF_stage/reg_bank/U1744  ( .A(\iRF_stage/reg_bank/n1701 ), .B(
        \iRF_stage/reg_bank/n1696 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1099 ) );
  MX4X1 \iRF_stage/reg_bank/U1749  ( .A(\iRF_stage/reg_bank/n1705 ), .B(
        \iRF_stage/reg_bank/n1703 ), .C(\iRF_stage/reg_bank/n1704 ), .D(
        \iRF_stage/reg_bank/n1702 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1706 ) );
  MX2X2 \iRF_stage/reg_bank/U1755  ( .A(\iRF_stage/reg_bank/n1711 ), .B(
        \iRF_stage/reg_bank/n1706 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1098 ) );
  MX4X1 \iRF_stage/reg_bank/U1760  ( .A(\iRF_stage/reg_bank/n1715 ), .B(
        \iRF_stage/reg_bank/n1713 ), .C(\iRF_stage/reg_bank/n1714 ), .D(
        \iRF_stage/reg_bank/n1712 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1716 ) );
  MX2X2 \iRF_stage/reg_bank/U1766  ( .A(\iRF_stage/reg_bank/n1721 ), .B(
        \iRF_stage/reg_bank/n1716 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1097 ) );
  MX4X1 \iRF_stage/reg_bank/U1771  ( .A(\iRF_stage/reg_bank/n1725 ), .B(
        \iRF_stage/reg_bank/n1723 ), .C(\iRF_stage/reg_bank/n1724 ), .D(
        \iRF_stage/reg_bank/n1722 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1726 ) );
  MX2X2 \iRF_stage/reg_bank/U1777  ( .A(\iRF_stage/reg_bank/n1731 ), .B(
        \iRF_stage/reg_bank/n1726 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1096 ) );
  MX4X1 \iRF_stage/reg_bank/U1782  ( .A(\iRF_stage/reg_bank/n1735 ), .B(
        \iRF_stage/reg_bank/n1733 ), .C(\iRF_stage/reg_bank/n1734 ), .D(
        \iRF_stage/reg_bank/n1732 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1736 ) );
  MX2X2 \iRF_stage/reg_bank/U1788  ( .A(\iRF_stage/reg_bank/n1741 ), .B(
        \iRF_stage/reg_bank/n1736 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1095 ) );
  MX4X1 \iRF_stage/reg_bank/U1793  ( .A(\iRF_stage/reg_bank/n1745 ), .B(
        \iRF_stage/reg_bank/n1743 ), .C(\iRF_stage/reg_bank/n1744 ), .D(
        \iRF_stage/reg_bank/n1742 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1746 ) );
  MX2X2 \iRF_stage/reg_bank/U1799  ( .A(\iRF_stage/reg_bank/n1751 ), .B(
        \iRF_stage/reg_bank/n1746 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1094 ) );
  MX4X1 \iRF_stage/reg_bank/U1804  ( .A(\iRF_stage/reg_bank/n1755 ), .B(
        \iRF_stage/reg_bank/n1753 ), .C(\iRF_stage/reg_bank/n1754 ), .D(
        \iRF_stage/reg_bank/n1752 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1756 ) );
  MX2X2 \iRF_stage/reg_bank/U1810  ( .A(\iRF_stage/reg_bank/n1761 ), .B(
        \iRF_stage/reg_bank/n1756 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1093 ) );
  MX4X1 \iRF_stage/reg_bank/U1815  ( .A(\iRF_stage/reg_bank/n1765 ), .B(
        \iRF_stage/reg_bank/n1763 ), .C(\iRF_stage/reg_bank/n1764 ), .D(
        \iRF_stage/reg_bank/n1762 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1766 ) );
  MX2X2 \iRF_stage/reg_bank/U1821  ( .A(\iRF_stage/reg_bank/n1771 ), .B(
        \iRF_stage/reg_bank/n1766 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1092 ) );
  MX4X1 \iRF_stage/reg_bank/U1826  ( .A(\iRF_stage/reg_bank/n1775 ), .B(
        \iRF_stage/reg_bank/n1773 ), .C(\iRF_stage/reg_bank/n1774 ), .D(
        \iRF_stage/reg_bank/n1772 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1776 ) );
  MX2X2 \iRF_stage/reg_bank/U1832  ( .A(\iRF_stage/reg_bank/n1781 ), .B(
        \iRF_stage/reg_bank/n1776 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1091 ) );
  MX4X1 \iRF_stage/reg_bank/U1837  ( .A(\iRF_stage/reg_bank/n1785 ), .B(
        \iRF_stage/reg_bank/n1783 ), .C(\iRF_stage/reg_bank/n1784 ), .D(
        \iRF_stage/reg_bank/n1782 ), .S0(\iRF_stage/reg_bank/N20 ), .S1(
        \iRF_stage/reg_bank/N19 ), .Y(\iRF_stage/reg_bank/n1786 ) );
  MX2X2 \iRF_stage/reg_bank/U1843  ( .A(\iRF_stage/reg_bank/n1791 ), .B(
        \iRF_stage/reg_bank/n1786 ), .S0(\iRF_stage/reg_bank/N21 ), .Y(
        \iRF_stage/reg_bank/N1090 ) );
  MX4XL \iRF_stage/reg_bank/U1265  ( .A(\iRF_stage/reg_bank/n1265 ), .B(
        \iRF_stage/reg_bank/n1263 ), .C(\iRF_stage/reg_bank/n1264 ), .D(
        \iRF_stage/reg_bank/n1262 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1266 ) );
  MX2X2 \iRF_stage/reg_bank/U1271  ( .A(\iRF_stage/reg_bank/n1271 ), .B(
        \iRF_stage/reg_bank/n1266 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1073 ) );
  MX4XL \iRF_stage/reg_bank/U1276  ( .A(\iRF_stage/reg_bank/n1275 ), .B(
        \iRF_stage/reg_bank/n1273 ), .C(\iRF_stage/reg_bank/n1274 ), .D(
        \iRF_stage/reg_bank/n1272 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1276 ) );
  MX2X2 \iRF_stage/reg_bank/U1282  ( .A(\iRF_stage/reg_bank/n1281 ), .B(
        \iRF_stage/reg_bank/n1276 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1072 ) );
  MX4X1 \iRF_stage/reg_bank/U1155  ( .A(\iRF_stage/reg_bank/n1165 ), .B(
        \iRF_stage/reg_bank/n1163 ), .C(\iRF_stage/reg_bank/n1164 ), .D(
        \iRF_stage/reg_bank/n1162 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1166 ) );
  MX2X2 \iRF_stage/reg_bank/U1161  ( .A(\iRF_stage/reg_bank/n1171 ), .B(
        \iRF_stage/reg_bank/n1166 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1083 ) );
  MX4X1 \iRF_stage/reg_bank/U1496  ( .A(\iRF_stage/reg_bank/n1475 ), .B(
        \iRF_stage/reg_bank/n1473 ), .C(\iRF_stage/reg_bank/n1474 ), .D(
        \iRF_stage/reg_bank/n1472 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1476 ) );
  MX2X2 \iRF_stage/reg_bank/U1502  ( .A(\iRF_stage/reg_bank/n1481 ), .B(
        \iRF_stage/reg_bank/n1476 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1052 ) );
  MX4X1 \iRF_stage/reg_bank/U1177  ( .A(\iRF_stage/reg_bank/n1185 ), .B(
        \iRF_stage/reg_bank/n1183 ), .C(\iRF_stage/reg_bank/n1184 ), .D(
        \iRF_stage/reg_bank/n1182 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1186 ) );
  MX2X2 \iRF_stage/reg_bank/U1183  ( .A(\iRF_stage/reg_bank/n1191 ), .B(
        \iRF_stage/reg_bank/n1186 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1081 ) );
  MX4X1 \iRF_stage/reg_bank/U1221  ( .A(\iRF_stage/reg_bank/n1225 ), .B(
        \iRF_stage/reg_bank/n1223 ), .C(\iRF_stage/reg_bank/n1224 ), .D(
        \iRF_stage/reg_bank/n1222 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1226 ) );
  MX2X2 \iRF_stage/reg_bank/U1227  ( .A(\iRF_stage/reg_bank/n1231 ), .B(
        \iRF_stage/reg_bank/n1226 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1077 ) );
  MX4X1 \iRF_stage/reg_bank/U1287  ( .A(\iRF_stage/reg_bank/n1285 ), .B(
        \iRF_stage/reg_bank/n1283 ), .C(\iRF_stage/reg_bank/n1284 ), .D(
        \iRF_stage/reg_bank/n1282 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1286 ) );
  MX2X2 \iRF_stage/reg_bank/U1293  ( .A(\iRF_stage/reg_bank/n1291 ), .B(
        \iRF_stage/reg_bank/n1286 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1071 ) );
  MX4X1 \iRF_stage/reg_bank/U1331  ( .A(\iRF_stage/reg_bank/n1325 ), .B(
        \iRF_stage/reg_bank/n1323 ), .C(\iRF_stage/reg_bank/n1324 ), .D(
        \iRF_stage/reg_bank/n1322 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1326 ) );
  MX2X2 \iRF_stage/reg_bank/U1337  ( .A(\iRF_stage/reg_bank/n1331 ), .B(
        \iRF_stage/reg_bank/n1326 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1067 ) );
  MX4X1 \iRF_stage/reg_bank/U1408  ( .A(\iRF_stage/reg_bank/n1395 ), .B(
        \iRF_stage/reg_bank/n1393 ), .C(\iRF_stage/reg_bank/n1394 ), .D(
        \iRF_stage/reg_bank/n1392 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1396 ) );
  MX2X2 \iRF_stage/reg_bank/U1414  ( .A(\iRF_stage/reg_bank/n1401 ), .B(
        \iRF_stage/reg_bank/n1396 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1060 ) );
  MX4X1 \iRF_stage/reg_bank/U1452  ( .A(\iRF_stage/reg_bank/n1435 ), .B(
        \iRF_stage/reg_bank/n1433 ), .C(\iRF_stage/reg_bank/n1434 ), .D(
        \iRF_stage/reg_bank/n1432 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1436 ) );
  MX2X2 \iRF_stage/reg_bank/U1458  ( .A(\iRF_stage/reg_bank/n1441 ), .B(
        \iRF_stage/reg_bank/n1436 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1056 ) );
  MX4X1 \iRF_stage/reg_bank/U1199  ( .A(\iRF_stage/reg_bank/n1205 ), .B(
        \iRF_stage/reg_bank/n1203 ), .C(\iRF_stage/reg_bank/n1204 ), .D(
        \iRF_stage/reg_bank/n1202 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1206 ) );
  MX2X2 \iRF_stage/reg_bank/U1205  ( .A(\iRF_stage/reg_bank/n1211 ), .B(
        \iRF_stage/reg_bank/n1206 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1079 ) );
  MX4X1 \iRF_stage/reg_bank/U1243  ( .A(\iRF_stage/reg_bank/n1245 ), .B(
        \iRF_stage/reg_bank/n1243 ), .C(\iRF_stage/reg_bank/n1244 ), .D(
        \iRF_stage/reg_bank/n1242 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1246 ) );
  MX2X2 \iRF_stage/reg_bank/U1249  ( .A(\iRF_stage/reg_bank/n1251 ), .B(
        \iRF_stage/reg_bank/n1246 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1075 ) );
  MX4X1 \iRF_stage/reg_bank/U1309  ( .A(\iRF_stage/reg_bank/n1305 ), .B(
        \iRF_stage/reg_bank/n1303 ), .C(\iRF_stage/reg_bank/n1304 ), .D(
        \iRF_stage/reg_bank/n1302 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1306 ) );
  MX2X2 \iRF_stage/reg_bank/U1315  ( .A(\iRF_stage/reg_bank/n1311 ), .B(
        \iRF_stage/reg_bank/n1306 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1069 ) );
  MX4X1 \iRF_stage/reg_bank/U1353  ( .A(\iRF_stage/reg_bank/n1345 ), .B(
        \iRF_stage/reg_bank/n1343 ), .C(\iRF_stage/reg_bank/n1344 ), .D(
        \iRF_stage/reg_bank/n1342 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1346 ) );
  MX2X2 \iRF_stage/reg_bank/U1359  ( .A(\iRF_stage/reg_bank/n1351 ), .B(
        \iRF_stage/reg_bank/n1346 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1065 ) );
  MX4X1 \iRF_stage/reg_bank/U1386  ( .A(\iRF_stage/reg_bank/n1375 ), .B(
        \iRF_stage/reg_bank/n1373 ), .C(\iRF_stage/reg_bank/n1374 ), .D(
        \iRF_stage/reg_bank/n1372 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1376 ) );
  MX2X2 \iRF_stage/reg_bank/U1392  ( .A(\iRF_stage/reg_bank/n1381 ), .B(
        \iRF_stage/reg_bank/n1376 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1062 ) );
  MX4X1 \iRF_stage/reg_bank/U1430  ( .A(\iRF_stage/reg_bank/n1415 ), .B(
        \iRF_stage/reg_bank/n1413 ), .C(\iRF_stage/reg_bank/n1414 ), .D(
        \iRF_stage/reg_bank/n1412 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1416 ) );
  MX2X2 \iRF_stage/reg_bank/U1436  ( .A(\iRF_stage/reg_bank/n1421 ), .B(
        \iRF_stage/reg_bank/n1416 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1058 ) );
  MX4X1 \iRF_stage/reg_bank/U1188  ( .A(\iRF_stage/reg_bank/n1195 ), .B(
        \iRF_stage/reg_bank/n1193 ), .C(\iRF_stage/reg_bank/n1194 ), .D(
        \iRF_stage/reg_bank/n1192 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1196 ) );
  MX2X2 \iRF_stage/reg_bank/U1194  ( .A(\iRF_stage/reg_bank/n1201 ), .B(
        \iRF_stage/reg_bank/n1196 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1080 ) );
  MX4X1 \iRF_stage/reg_bank/U1232  ( .A(\iRF_stage/reg_bank/n1235 ), .B(
        \iRF_stage/reg_bank/n1233 ), .C(\iRF_stage/reg_bank/n1234 ), .D(
        \iRF_stage/reg_bank/n1232 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1236 ) );
  MX2X2 \iRF_stage/reg_bank/U1238  ( .A(\iRF_stage/reg_bank/n1241 ), .B(
        \iRF_stage/reg_bank/n1236 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1076 ) );
  MX4X1 \iRF_stage/reg_bank/U1298  ( .A(\iRF_stage/reg_bank/n1295 ), .B(
        \iRF_stage/reg_bank/n1293 ), .C(\iRF_stage/reg_bank/n1294 ), .D(
        \iRF_stage/reg_bank/n1292 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1296 ) );
  MX2X2 \iRF_stage/reg_bank/U1304  ( .A(\iRF_stage/reg_bank/n1301 ), .B(
        \iRF_stage/reg_bank/n1296 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1070 ) );
  MX4X1 \iRF_stage/reg_bank/U1342  ( .A(\iRF_stage/reg_bank/n1335 ), .B(
        \iRF_stage/reg_bank/n1333 ), .C(\iRF_stage/reg_bank/n1334 ), .D(
        \iRF_stage/reg_bank/n1332 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1336 ) );
  MX2X2 \iRF_stage/reg_bank/U1348  ( .A(\iRF_stage/reg_bank/n1341 ), .B(
        \iRF_stage/reg_bank/n1336 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1066 ) );
  MX4X1 \iRF_stage/reg_bank/U1375  ( .A(\iRF_stage/reg_bank/n1365 ), .B(
        \iRF_stage/reg_bank/n1363 ), .C(\iRF_stage/reg_bank/n1364 ), .D(
        \iRF_stage/reg_bank/n1362 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1366 ) );
  MX2X2 \iRF_stage/reg_bank/U1381  ( .A(\iRF_stage/reg_bank/n1371 ), .B(
        \iRF_stage/reg_bank/n1366 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1063 ) );
  MX4X1 \iRF_stage/reg_bank/U1419  ( .A(\iRF_stage/reg_bank/n1405 ), .B(
        \iRF_stage/reg_bank/n1403 ), .C(\iRF_stage/reg_bank/n1404 ), .D(
        \iRF_stage/reg_bank/n1402 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1406 ) );
  MX2X2 \iRF_stage/reg_bank/U1425  ( .A(\iRF_stage/reg_bank/n1411 ), .B(
        \iRF_stage/reg_bank/n1406 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1059 ) );
  MX4X1 \iRF_stage/reg_bank/U1210  ( .A(\iRF_stage/reg_bank/n1215 ), .B(
        \iRF_stage/reg_bank/n1213 ), .C(\iRF_stage/reg_bank/n1214 ), .D(
        \iRF_stage/reg_bank/n1212 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1216 ) );
  MX2X2 \iRF_stage/reg_bank/U1216  ( .A(\iRF_stage/reg_bank/n1221 ), .B(
        \iRF_stage/reg_bank/n1216 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1078 ) );
  MX4X1 \iRF_stage/reg_bank/U1254  ( .A(\iRF_stage/reg_bank/n1255 ), .B(
        \iRF_stage/reg_bank/n1253 ), .C(\iRF_stage/reg_bank/n1254 ), .D(
        \iRF_stage/reg_bank/n1252 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1256 ) );
  MX2X2 \iRF_stage/reg_bank/U1260  ( .A(\iRF_stage/reg_bank/n1261 ), .B(
        \iRF_stage/reg_bank/n1256 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1074 ) );
  MX4X1 \iRF_stage/reg_bank/U1320  ( .A(\iRF_stage/reg_bank/n1315 ), .B(
        \iRF_stage/reg_bank/n1313 ), .C(\iRF_stage/reg_bank/n1314 ), .D(
        \iRF_stage/reg_bank/n1312 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1316 ) );
  MX2X2 \iRF_stage/reg_bank/U1326  ( .A(\iRF_stage/reg_bank/n1321 ), .B(
        \iRF_stage/reg_bank/n1316 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1068 ) );
  MX4X1 \iRF_stage/reg_bank/U1364  ( .A(\iRF_stage/reg_bank/n1355 ), .B(
        \iRF_stage/reg_bank/n1353 ), .C(\iRF_stage/reg_bank/n1354 ), .D(
        \iRF_stage/reg_bank/n1352 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1356 ) );
  MX2X2 \iRF_stage/reg_bank/U1370  ( .A(\iRF_stage/reg_bank/n1361 ), .B(
        \iRF_stage/reg_bank/n1356 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1064 ) );
  MX4X1 \iRF_stage/reg_bank/U1397  ( .A(\iRF_stage/reg_bank/n1385 ), .B(
        \iRF_stage/reg_bank/n1383 ), .C(\iRF_stage/reg_bank/n1384 ), .D(
        \iRF_stage/reg_bank/n1382 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1386 ) );
  MX2X2 \iRF_stage/reg_bank/U1403  ( .A(\iRF_stage/reg_bank/n1391 ), .B(
        \iRF_stage/reg_bank/n1386 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1061 ) );
  MX4X1 \iRF_stage/reg_bank/U1441  ( .A(\iRF_stage/reg_bank/n1425 ), .B(
        \iRF_stage/reg_bank/n1423 ), .C(\iRF_stage/reg_bank/n1424 ), .D(
        \iRF_stage/reg_bank/n1422 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1426 ) );
  MX2X2 \iRF_stage/reg_bank/U1447  ( .A(\iRF_stage/reg_bank/n1431 ), .B(
        \iRF_stage/reg_bank/n1426 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1057 ) );
  MX4X1 \iRF_stage/reg_bank/U1166  ( .A(\iRF_stage/reg_bank/n1175 ), .B(
        \iRF_stage/reg_bank/n1173 ), .C(\iRF_stage/reg_bank/n1174 ), .D(
        \iRF_stage/reg_bank/n1172 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1176 ) );
  MX2X2 \iRF_stage/reg_bank/U1172  ( .A(\iRF_stage/reg_bank/n1181 ), .B(
        \iRF_stage/reg_bank/n1176 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1082 ) );
  MX4X1 \iRF_stage/reg_bank/U1485  ( .A(\iRF_stage/reg_bank/n1465 ), .B(
        \iRF_stage/reg_bank/n1463 ), .C(\iRF_stage/reg_bank/n1464 ), .D(
        \iRF_stage/reg_bank/n1462 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1466 ) );
  MX2X2 \iRF_stage/reg_bank/U1491  ( .A(\iRF_stage/reg_bank/n1471 ), .B(
        \iRF_stage/reg_bank/n1466 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1053 ) );
  MX4X1 \iRF_stage/reg_bank/U1474  ( .A(\iRF_stage/reg_bank/n1455 ), .B(
        \iRF_stage/reg_bank/n1453 ), .C(\iRF_stage/reg_bank/n1454 ), .D(
        \iRF_stage/reg_bank/n1452 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1456 ) );
  MX2X2 \iRF_stage/reg_bank/U1480  ( .A(\iRF_stage/reg_bank/n1461 ), .B(
        \iRF_stage/reg_bank/n1456 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1054 ) );
  MX4X1 \iRF_stage/reg_bank/U1463  ( .A(\iRF_stage/reg_bank/n1445 ), .B(
        \iRF_stage/reg_bank/n1443 ), .C(\iRF_stage/reg_bank/n1444 ), .D(
        \iRF_stage/reg_bank/n1442 ), .S0(\iRF_stage/reg_bank/N15 ), .S1(
        \iRF_stage/reg_bank/N14 ), .Y(\iRF_stage/reg_bank/n1446 ) );
  MX2X2 \iRF_stage/reg_bank/U1469  ( .A(\iRF_stage/reg_bank/n1451 ), .B(
        \iRF_stage/reg_bank/n1446 ), .S0(\iRF_stage/reg_bank/N16 ), .Y(
        \iRF_stage/reg_bank/N1055 ) );
  EDFFTRX1 \decoder_pipe/pipereg/U1/muxb_ctl_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2094[0] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5483[0] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U1/muxb_ctl_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2094[1] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5483[1] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U26/alu_func_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2040[0] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5674[0] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U26/alu_func_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2040[1] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5674[1] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U26/alu_func_o_reg_2_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2040[2] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5674[2] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U26/alu_func_o_reg_3_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2040[3] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5674[3] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U26/alu_func_o_reg_4_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2040[4] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5674[4] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U3/dmem_ctl_o_reg_0_  ( .RN(n1933), .D(n1928), 
        .E(n1936), .CK(clk), .Q(\decoder_pipe/pipereg/BUS5666[0] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U3/dmem_ctl_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2064[1] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5666[1] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U3/dmem_ctl_o_reg_2_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2064[2] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5666[2] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U3/dmem_ctl_o_reg_3_  ( .RN(n1933), .D(n1931), 
        .E(n1936), .CK(clk), .Q(\decoder_pipe/pipereg/BUS5666[3] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U7/muxa_ctl_o_reg_0_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2086[0] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5008[0] ) );
  EDFFTRX1 \decoder_pipe/pipereg/U7/muxa_ctl_o_reg_1_  ( .RN(n1933), .D(
        \decoder_pipe/BUS2086[1] ), .E(n1936), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5008[1] ) );
  DFFHQX1 \rnd_pass0/r5_o_reg_0_  ( .D(BUS775[0]), .CK(clk), .Q(BUS1726[0]) );
  DFFHQX1 \rnd_pass0/r5_o_reg_1_  ( .D(BUS775[1]), .CK(clk), .Q(BUS1726[1]) );
  DFFHQX1 \rnd_pass0/r5_o_reg_2_  ( .D(BUS775[2]), .CK(clk), .Q(BUS1726[2]) );
  DFFHQX1 \rnd_pass0/r5_o_reg_3_  ( .D(BUS775[3]), .CK(clk), .Q(BUS1726[3]) );
  DFFHQX1 \rnd_pass0/r5_o_reg_4_  ( .D(BUS775[4]), .CK(clk), .Q(BUS1726[4]) );
  XOR3X2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_31  ( .A(
        \iexec_stage/BUS476[31] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[31] ), .C(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[31] ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/N143 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_2  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_2 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_2 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[2] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[3] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N178 ) );
  ADDFXL \iexec_stage/MIPS_alu/mips_alu/r92/U1_2  ( .A(\iexec_stage/BUS476[2] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[2] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[2] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[3] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N114 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_3  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_3 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_3 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[3] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[4] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N179 ) );
  ADDFXL \iexec_stage/MIPS_alu/mips_alu/r92/U1_3  ( .A(\iexec_stage/BUS476[3] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[3] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[3] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[4] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N115 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_10  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_10 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_10 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[10] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[11] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N186 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_10  ( .A(
        \iexec_stage/BUS476[10] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[10] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[10] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[11] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N122 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_16  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_16 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_16 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[16] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[17] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N192 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_16  ( .A(
        \iexec_stage/BUS476[16] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[16] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[16] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[17] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N128 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_17  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_17 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_17 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[17] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[18] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N193 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_17  ( .A(
        \iexec_stage/BUS476[17] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[17] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[17] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[18] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N129 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_18  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_18 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_18 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[18] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[19] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N194 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_18  ( .A(
        \iexec_stage/BUS476[18] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[18] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[18] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[19] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N130 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_19  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_19 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_19 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[19] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[20] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N195 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_19  ( .A(
        \iexec_stage/BUS476[19] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[19] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[19] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[20] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N131 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_20  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_20 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_20 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[20] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[21] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N196 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_20  ( .A(
        \iexec_stage/BUS476[20] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[20] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[20] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[21] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N132 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_21  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_21 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_21 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[21] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[22] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N197 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_21  ( .A(
        \iexec_stage/BUS476[21] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[21] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[21] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[22] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N133 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_22  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_22 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_22 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[22] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[23] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N198 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_22  ( .A(
        \iexec_stage/BUS476[22] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[22] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[22] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[23] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N134 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_23  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_23 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_23 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[23] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[24] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N199 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_23  ( .A(
        \iexec_stage/BUS476[23] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[23] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[23] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[24] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N135 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_24  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_24 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_24 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[24] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[25] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N200 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_24  ( .A(
        \iexec_stage/BUS476[24] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[24] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[24] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[25] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N136 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_25  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_25 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_25 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[25] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[26] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N201 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_26  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_26 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_26 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[26] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[27] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N202 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_27  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_27 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_27 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[27] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[28] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N203 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_28  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_28 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_28 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[28] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[29] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N204 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_30  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_30 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_30 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[30] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[31] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N206 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_30  ( .A(
        \iexec_stage/BUS476[30] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[30] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[30] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[31] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N142 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_31  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_32 ), .B(n1879), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[31] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[32] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N207 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_9  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_9 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_9 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[9] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[10] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N185 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_15  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_15 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_15 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[15] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[16] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N191 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_29  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_29 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_29 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[29] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[30] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N205 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_8  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_8 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_8 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[8] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[9] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N184 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_14  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_14 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_14 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[14] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[15] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N190 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_7  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_7 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_7 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[7] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[8] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N183 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_9  ( .A(\iexec_stage/BUS476[9] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[9] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[9] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[10] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N121 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_13  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_13 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_13 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[13] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[14] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N189 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_15  ( .A(
        \iexec_stage/BUS476[15] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[15] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[15] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[16] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N127 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_29  ( .A(
        \iexec_stage/BUS476[29] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[29] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[29] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[30] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N141 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_6  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_6 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_6 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[6] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[7] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N182 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_8  ( .A(\iexec_stage/BUS476[8] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[8] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[8] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[9] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N120 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_12  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_12 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_12 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[12] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[13] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N188 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_14  ( .A(
        \iexec_stage/BUS476[14] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[14] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[14] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[15] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N126 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_28  ( .A(
        \iexec_stage/BUS476[28] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[28] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[28] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[29] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N140 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_5  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_5 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_5 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[5] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[6] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N181 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_7  ( .A(\iexec_stage/BUS476[7] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[7] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[7] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[8] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N119 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_11  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_11 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_11 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[11] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[12] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N187 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_13  ( .A(
        \iexec_stage/BUS476[13] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[13] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[13] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[14] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N125 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_27  ( .A(
        \iexec_stage/BUS476[27] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[27] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[27] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[28] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N139 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_4  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_4 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_4 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[4] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[5] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N180 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_6  ( .A(\iexec_stage/BUS476[6] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[6] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[6] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[7] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N118 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_12  ( .A(
        \iexec_stage/BUS476[12] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[12] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[12] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[13] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N124 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_26  ( .A(
        \iexec_stage/BUS476[26] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[26] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[26] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[27] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N138 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_5  ( .A(\iexec_stage/BUS476[5] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[5] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[5] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[6] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N117 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_11  ( .A(
        \iexec_stage/BUS476[11] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[11] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[11] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[12] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N123 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r92/U1_25  ( .A(
        \iexec_stage/BUS476[25] ), .B(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[25] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[25] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[26] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N137 ) );
  ADDFXL \iexec_stage/MIPS_alu/mips_alu/r92/U1_4  ( .A(\iexec_stage/BUS476[4] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[4] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[4] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[5] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N116 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_1  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_1 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_1 ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[1] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[2] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N177 ) );
  ADDFXL \iexec_stage/MIPS_alu/mips_alu/r92/U1_1  ( .A(\iexec_stage/BUS476[1] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[1] ), .CI(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[1] ), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[2] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N113 ) );
  ADDFX2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_0  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_0 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_0 ), .CI(n1938), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[1] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N176 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U462  ( .A(n116), .B(n119), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N202 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U461  ( .A(n115), .B(n118), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N203 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U460  ( .A(n114), .B(n117), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N204 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U428  ( .A(n87), .B(n105), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N242 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U427  ( .A(n86), .B(n103), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N243 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U426  ( .A(n85), .B(n93), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N244 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U453  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n407 ), .B(n1884), .S0(
        \iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n408 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U454  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n408 ), .B(n111), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n409 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U455  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n409 ), .B(n114), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N208 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U458  ( .A(n107), .B(n1888), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n411 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U459  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n411 ), .B(n113), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N205 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U424  ( .A(n105), .B(n102), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N246 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U423  ( .A(n103), .B(n100), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N247 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U422  ( .A(n93), .B(n90), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N248 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U419  ( .A(n102), .B(n98), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N250 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U438  ( .A(n99), .B(n95), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N219 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U416  ( .A(n1890), .B(
        \iexec_stage/BUS468[31] ), .S0(\iexec_stage/BUS476[4] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n398 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U417  ( .A(n90), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n398 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N252 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U412  ( .A(n124), .B(
        \iexec_stage/BUS468[31] ), .S0(\iexec_stage/BUS476[4] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n396 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U413  ( .A(n98), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n396 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N254 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U410  ( .A(n123), .B(
        \iexec_stage/BUS468[31] ), .S0(\iexec_stage/BUS476[4] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n395 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U411  ( .A(n96), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n395 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N255 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U678  ( .A(n1914), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n600 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n601 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U679  ( .A(n110), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n601 ), .S0(\iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n427 ) );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U482  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n427 ), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n426 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U483  ( .A(n122), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n426 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N193 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U673  ( .A(n1908), .B(n108), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n419 )
         );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U474  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n419 ), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n418 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U475  ( .A(n121), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n418 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N196 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U473  ( .A(n120), .B(n122), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N197 )
         );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U469  ( .A(n1910), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n415 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U470  ( .A(n1904), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n415 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n416 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U471  ( .A(n82), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n416 ), .S0(\iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n417 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U472  ( .A(n119), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n417 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N198 ) );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U465  ( .A(n1907), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n412 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U466  ( .A(n1902), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n412 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n413 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U467  ( .A(n1900), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n413 ), .S0(\iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n414 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U468  ( .A(n118), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n414 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N199 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U464  ( .A(n117), .B(n121), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N200 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U463  ( .A(n113), .B(n120), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N201 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U456  ( .A(n112), .B(n107), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n410 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U457  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n410 ), .B(n116), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N206 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U444  ( .A(n106), .B(n101), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N214 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U443  ( .A(n104), .B(n99), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N215 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U442  ( .A(n94), .B(n89), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N216 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U439  ( .A(n101), .B(n97), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N218 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U418  ( .A(n100), .B(n96), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N251 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U437  ( .A(n89), .B(n88), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N220 )
         );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U433  ( .A(n124), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n402 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U434  ( .A(n97), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n402 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N222 ) );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U431  ( .A(n123), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n401 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U432  ( .A(n95), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n401 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N223 ) );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U429  ( .A(n1882), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n400 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U430  ( .A(n88), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n400 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N224 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U402  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n387 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n384 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n386 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U401  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n384 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n385 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n383 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U403  ( .A(\iexec_stage/BUS476[0] ), 
        .B(n1881), .Y(\iexec_stage/MIPS_alu/mips_shifter/n388 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U529  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n457 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n387 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n458 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U449  ( .A(n111), .B(n112), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n405 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U574  ( .A(n1926), .B(n1925), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n503 )
         );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U404  ( .A(\iexec_stage/BUS476[1] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n388 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n389 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U445  ( .A(n84), .B(n92), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N213 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U425  ( .A(n84), .B(n91), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N245 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U420  ( .A(n1894), .B(
        \iexec_stage/BUS468[31] ), .S0(\iexec_stage/BUS476[4] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n399 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U421  ( .A(n1880), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n399 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N249 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U414  ( .A(n1887), .B(
        \iexec_stage/BUS468[31] ), .S0(\iexec_stage/BUS476[4] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n397 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U415  ( .A(n91), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n397 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N253 ) );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U440  ( .A(n1894), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n404 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U441  ( .A(n1880), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n404 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N217 ) );
  AND2X1 \iexec_stage/MIPS_alu/mips_shifter/U435  ( .A(n1887), .B(n1923), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n403 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U436  ( .A(n92), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n403 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N221 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U488  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1909), .Y(\iexec_stage/MIPS_alu/mips_shifter/n434 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U489  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1911), .Y(\iexec_stage/MIPS_alu/mips_shifter/n435 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U408  ( .A(n1890), .B(n1882), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n394 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U409  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n394 ), .B(\iexec_stage/BUS468[31] ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N256 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U677  ( .A(\iexec_stage/BUS468[9] ), 
        .B(\iexec_stage/BUS468[1] ), .S0(\iexec_stage/BUS476[3] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n600 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U578  ( .A(n1927), .B(n1926), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n507 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U579  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n507 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n499 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n508 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U580  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n508 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n492 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n509 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U581  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n509 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n386 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n510 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U570  ( .A(n1925), .B(n1924), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n499 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U562  ( .A(n1922), .B(n1921), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n491 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U554  ( .A(n1920), .B(n1919), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n483 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U511  ( .A(n1906), .B(n1903), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n444 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U506  ( .A(n1901), .B(n1899), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n369 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U505  ( .A(n1898), .B(n1897), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n370 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U508  ( .A(n1896), .B(n1895), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n366 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U519  ( .A(n1912), .B(n1911), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n451 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U499  ( .A(n1909), .B(n1906), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n438 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U558  ( .A(n1921), .B(n1920), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n487 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U550  ( .A(n1919), .B(n1918), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n479 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U492  ( .A(n1897), .B(n1896), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n374 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U496  ( .A(n1895), .B(n1893), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n375 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U566  ( .A(n1924), .B(n1922), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n495 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U498  ( .A(n1903), .B(n1901), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n377 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U493  ( .A(n1899), .B(n1898), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n378 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U542  ( .A(n1917), .B(n1916), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n471 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U532  ( .A(n1915), .B(n1913), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n461 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U495  ( .A(n1892), .B(n1891), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n436 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U491  ( .A(n1889), .B(n1886), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n360 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U512  ( .A(n1911), .B(n1909), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n445 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U546  ( .A(n1918), .B(n1917), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n475 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U507  ( .A(n1893), .B(n1892), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n367 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U537  ( .A(n1916), .B(n1915), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n466 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U527  ( .A(n1913), .B(n1912), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n456 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U503  ( .A(n1891), .B(n1889), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n441 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U502  ( .A(n1886), .B(n1885), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n382 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U661  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n581 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n589 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n590 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U407  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n390 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n393 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n392 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U392  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n363 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n359 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n362 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U485  ( .A(n1915), .B(n1924), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n431 )
         );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U667  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1920), .Y(\iexec_stage/MIPS_alu/mips_shifter/n595 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U668  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n435 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n595 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n596 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U669  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n589 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n596 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n597 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U633  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n550 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n538 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n562 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U501  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n439 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n437 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n440 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U623  ( .A(n1885), .B(n1912), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n552 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U624  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n552 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n551 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n553 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U405  ( .A(n1909), .B(n1919), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n390 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U406  ( .A(n1911), .B(n1920), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n391 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U605  ( .A(n1895), .B(n1919), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n534 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U516  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n436 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n360 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n380 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U504  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n441 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n382 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n372 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U523  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n367 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n441 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n385 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U547  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n475 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n466 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n476 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U657  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n577 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n585 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n586 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U653  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n573 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n581 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n582 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U649  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n569 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n577 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n578 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U645  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n564 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n573 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n574 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U610  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n538 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n535 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n539 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U617  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n545 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n542 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n546 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U563  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n491 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n483 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n492 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U526  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n444 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n369 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n387 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U524  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n370 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n366 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n384 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U500  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n438 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n377 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n439 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U533  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n461 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n451 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n462 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U494  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n378 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n374 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n363 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U636  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n542 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n564 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n565 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U641  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n535 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n569 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n570 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U528  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n456 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n445 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n457 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U651  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1916), .Y(\iexec_stage/MIPS_alu/mips_shifter/n580 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U652  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n543 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n580 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n581 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U647  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1915), .Y(\iexec_stage/MIPS_alu/mips_shifter/n576 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U648  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n548 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n576 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n577 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U643  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1913), .Y(\iexec_stage/MIPS_alu/mips_shifter/n572 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U644  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n555 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n572 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n573 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U672  ( .A(n1913), .B(n1922), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n429 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U666  ( .A(n1912), .B(n1921), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n393 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U612  ( .A(n1893), .B(n1918), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n541 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U613  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n541 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n540 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n542 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U635  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n558 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n435 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n564 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U606  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n534 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n434 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n535 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U639  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1912), .Y(\iexec_stage/MIPS_alu/mips_shifter/n568 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U640  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n551 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n568 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n569 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U620  ( .A(n1889), .B(n1915), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n549 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U621  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n549 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n548 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n550 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U608  ( .A(n1892), .B(n1917), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n537 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U609  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n537 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n536 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n538 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U627  ( .A(n1886), .B(n1913), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n556 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U628  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n556 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n555 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n557 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U615  ( .A(n1891), .B(n1916), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n544 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U616  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n544 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n543 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n545 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U520  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n451 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n438 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n452 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U513  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n445 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n444 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n446 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U589  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n361 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n388 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n518 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U590  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n452 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n518 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n519 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U518  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n361 ), .B(n1881), .S0(
        \iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n450 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U521  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n452 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n450 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n453 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U585  ( .A(\iexec_stage/BUS476[1] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n364 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n514 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U586  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n446 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n514 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n515 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U510  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n364 ), .B(n1881), .S0(
        \iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n443 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U514  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n446 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n443 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n447 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U629  ( .A(n1896), .B(n1920), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n558 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U611  ( .A(n1906), .B(n1927), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n540 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U622  ( .A(n1897), .B(n1921), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n551 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U619  ( .A(n1899), .B(n1924), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n548 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U607  ( .A(n1903), .B(n1926), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n536 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U626  ( .A(n1898), .B(n1922), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n555 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U614  ( .A(n1901), .B(n1925), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n543 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U551  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n479 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n471 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n480 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U552  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n480 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n439 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n481 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U534  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n462 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n363 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n463 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U393  ( .A(n1883), .B(n1881), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n364 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U559  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n487 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n479 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n488 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U560  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n488 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n373 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n489 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U555  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n483 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n475 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n484 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U556  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n484 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n365 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n485 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U490  ( .A(n1885), .B(n1883), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n361 )
         );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U659  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1918), .Y(\iexec_stage/MIPS_alu/mips_shifter/n588 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U660  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n540 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n588 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n589 ) );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U655  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1917), .Y(\iexec_stage/MIPS_alu/mips_shifter/n584 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U656  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n536 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n584 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n585 ) );
  MX4XL \iexec_stage/MIPS_alu/mips_shifter/U548  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n476 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n385 ), .C(
        \iexec_stage/MIPS_alu/mips_shifter/n457 ), .D(
        \iexec_stage/MIPS_alu/mips_shifter/n381 ), .S0(\iexec_stage/BUS476[4] ), .S1(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n477 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U397  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n374 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n375 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n373 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U394  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n366 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n367 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n365 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U391  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n360 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n361 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n359 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U400  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n382 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n364 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n381 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U497  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n375 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n436 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n437 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U543  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n471 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n461 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n472 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U544  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n472 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n380 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n473 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U538  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n466 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n456 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n467 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U539  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n467 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n372 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n468 ) );
  ADDFXL \iexec_stage/MIPS_alu/mips_alu/r92/U1_0  ( .A(\iexec_stage/BUS476[0] ), .B(\iexec_stage/MIPS_alu/mips_alu/r92/B_AS[0] ), .CI(n78), .CO(
        \iexec_stage/MIPS_alu/mips_alu/r92/carry[1] ), .S(
        \iexec_stage/MIPS_alu/mips_alu/N112 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U398  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n377 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n378 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n376 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U395  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n369 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n370 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n368 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U447  ( .A(n86), .B(n104), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N211 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U446  ( .A(n85), .B(n94), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N212 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U450  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n405 ), .B(n115), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N207 )
         );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U582  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n510 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n477 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n511 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U448  ( .A(n87), .B(n106), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/N210 )
         );
  XOR3X2 \iexec_stage/MIPS_alu/mips_alu/r86/U1_32  ( .A(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_32 ), .B(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_32 ), .C(
        \iexec_stage/MIPS_alu/mips_alu/r86/carry[32] ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/N370 ) );
  DFFHQX1 \cop_data_reg/r32_o_reg_0_  ( .D(dout[0]), .CK(clk), .Q(
        cop_data_o[0]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_1_  ( .D(dout[1]), .CK(clk), .Q(
        cop_data_o[1]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_2_  ( .D(dout[2]), .CK(clk), .Q(
        cop_data_o[2]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_3_  ( .D(dout[3]), .CK(clk), .Q(
        cop_data_o[3]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_4_  ( .D(dout[4]), .CK(clk), .Q(
        cop_data_o[4]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_5_  ( .D(dout[5]), .CK(clk), .Q(
        cop_data_o[5]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_6_  ( .D(dout[6]), .CK(clk), .Q(
        cop_data_o[6]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_7_  ( .D(dout[7]), .CK(clk), .Q(
        cop_data_o[7]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_8_  ( .D(BUS9884[8]), .CK(clk), .Q(
        cop_data_o[8]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_9_  ( .D(BUS9884[9]), .CK(clk), .Q(
        cop_data_o[9]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_10_  ( .D(BUS9884[10]), .CK(clk), .Q(
        cop_data_o[10]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_11_  ( .D(BUS9884[11]), .CK(clk), .Q(
        cop_data_o[11]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_12_  ( .D(BUS9884[12]), .CK(clk), .Q(
        cop_data_o[12]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_13_  ( .D(BUS9884[13]), .CK(clk), .Q(
        cop_data_o[13]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_14_  ( .D(BUS9884[14]), .CK(clk), .Q(
        cop_data_o[14]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_15_  ( .D(BUS9884[15]), .CK(clk), .Q(
        cop_data_o[15]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_16_  ( .D(BUS9884[16]), .CK(clk), .Q(
        cop_data_o[16]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_17_  ( .D(BUS9884[17]), .CK(clk), .Q(
        cop_data_o[17]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_18_  ( .D(BUS9884[18]), .CK(clk), .Q(
        cop_data_o[18]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_19_  ( .D(BUS9884[19]), .CK(clk), .Q(
        cop_data_o[19]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_20_  ( .D(BUS9884[20]), .CK(clk), .Q(
        cop_data_o[20]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_21_  ( .D(BUS9884[21]), .CK(clk), .Q(
        cop_data_o[21]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_22_  ( .D(BUS9884[22]), .CK(clk), .Q(
        cop_data_o[22]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_23_  ( .D(BUS9884[23]), .CK(clk), .Q(
        cop_data_o[23]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_24_  ( .D(BUS9884[24]), .CK(clk), .Q(
        cop_data_o[24]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_25_  ( .D(BUS9884[25]), .CK(clk), .Q(
        cop_data_o[25]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_26_  ( .D(BUS9884[26]), .CK(clk), .Q(
        cop_data_o[26]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_27_  ( .D(BUS9884[27]), .CK(clk), .Q(
        cop_data_o[27]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_28_  ( .D(BUS9884[28]), .CK(clk), .Q(
        cop_data_o[28]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_29_  ( .D(BUS9884[29]), .CK(clk), .Q(
        cop_data_o[29]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_30_  ( .D(BUS9884[30]), .CK(clk), .Q(
        cop_data_o[30]) );
  DFFHQX1 \cop_data_reg/r32_o_reg_31_  ( .D(BUS9884[31]), .CK(clk), .Q(
        cop_data_o[31]) );
  DFFTRX1 \decoder_pipe/pipereg/U13/wb_mux_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5651[0] ), .RN(n1934), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5690[0] ) );
  DFFTRX1 \decoder_pipe/pipereg/U19/wb_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5639[0] ), .RN(n1934), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5682[0] ) );
  DFFTRX1 \decoder_pipe/pipereg/U24/alu_we_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS4987[0] ), .RN(n1934), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS7299[0] ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U575  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n503 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n495 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n504 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U571  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n499 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n491 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n500 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U567  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n495 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n487 ), .S0(\iexec_stage/BUS476[1] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n496 ) );
  MX2X1 \iexec_stage/MIPS_alu/mips_shifter/U630  ( .A(n1883), .B(n1911), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n559 )
         );
  OR2XL \iexec_stage/MIPS_alu/mips_shifter/U663  ( .A(\iexec_stage/BUS476[4] ), 
        .B(n1919), .Y(\iexec_stage/MIPS_alu/mips_shifter/n592 ) );
  DFFHQX1 \decoder_pipe/pipereg/U9/dmem_ctl_o_reg_0_  ( .D(BUS5985[0]), .CK(
        clk), .Q(cop_mem_ctl_o[0]) );
  DFFHQX1 \decoder_pipe/pipereg/U9/dmem_ctl_o_reg_1_  ( .D(BUS5985[1]), .CK(
        clk), .Q(cop_mem_ctl_o[1]) );
  DFFHQX1 \decoder_pipe/pipereg/U9/dmem_ctl_o_reg_2_  ( .D(BUS5985[2]), .CK(
        clk), .Q(cop_mem_ctl_o[2]) );
  DFFHQX1 \decoder_pipe/pipereg/U9/dmem_ctl_o_reg_3_  ( .D(BUS5985[3]), .CK(
        clk), .Q(cop_mem_ctl_o[3]) );
  DFFHQX1 \decoder_pipe/pipereg/U21/wb_mux_ctl_o_reg_0_  ( .D(
        \decoder_pipe/pipereg/BUS5690[0] ), .CK(clk), .Q(
        \decoder_pipe/pipereg/BUS5790[0] ) );
  EDFFX2 \iRF_stage/reg_bank/r_rdaddress_b_reg_2_  ( .D(\iRF_stage/BUS3236[2] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N19 ), .QN(n341) );
  EDFFX2 \iRF_stage/reg_bank/r_rdaddress_a_reg_2_  ( .D(\iRF_stage/BUS3237[2] ), .E(n1936), .CK(clk), .Q(\iRF_stage/reg_bank/N14 ), .QN(n336) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U576  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n504 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n376 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n505 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U572  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n500 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n368 ), .S0(\iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n501 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U601  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n437 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n389 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n530 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U568  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n496 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n462 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n497 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U676  ( .A(n109), .B(n110), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n425 )
         );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U674  ( .A(n108), .B(n109), .S0(
        \iexec_stage/BUS476[0] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n422 )
         );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U549  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n437 ), .B(n1881), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n478 )
         );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U593  ( .A(\iexec_stage/BUS476[2] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n381 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n522 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U564  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n492 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n476 ), .S0(\iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n493 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U525  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n381 ), .B(n1881), .S0(
        \iexec_stage/BUS476[2] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n455 )
         );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U541  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n376 ), .B(n1881), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n470 )
         );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U599  ( .A(\iexec_stage/BUS476[4] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n376 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n528 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U536  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n368 ), .B(n1881), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n465 )
         );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U597  ( .A(\iexec_stage/BUS476[4] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n368 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n526 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U531  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n359 ), .B(n1881), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n460 )
         );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U595  ( .A(\iexec_stage/BUS476[3] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n359 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n524 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U517  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n373 ), .B(n1881), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n449 )
         );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U591  ( .A(\iexec_stage/BUS476[4] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n373 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n520 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U509  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n365 ), .B(n1881), .S0(
        \iexec_stage/BUS476[4] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n442 )
         );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U587  ( .A(\iexec_stage/BUS476[4] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n365 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n516 ) );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U583  ( .A(\iexec_stage/BUS476[3] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n389 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n512 ) );
  OR2X1 \iexec_stage/MIPS_alu/mips_shifter/U670  ( .A(\iexec_stage/BUS476[4] ), 
        .B(\iexec_stage/MIPS_alu/mips_shifter/n392 ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/n598 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U675  ( .A(n1916), .B(n1925), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n430 )
         );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U664  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n434 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n592 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n593 ) );
  MX2X2 \iexec_stage/MIPS_alu/mips_shifter/U631  ( .A(
        \iexec_stage/MIPS_alu/mips_shifter/n559 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n558 ), .S0(\iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n560 ) );
  OR4X2 U3 ( .A(n36), .B(n287), .C(n288), .D(n289), .Y(n1) );
  NAND2X2 U4 ( .A(n1547), .B(n1548), .Y(\iexec_stage/BUS476[1] ) );
  NAND2X2 U5 ( .A(n1545), .B(n1546), .Y(\iexec_stage/BUS476[3] ) );
  NAND2X2 U6 ( .A(n1551), .B(n1552), .Y(\iexec_stage/BUS476[4] ) );
  INVX2 U7 ( .A(n1), .Y(n78) );
  NAND2X2 U8 ( .A(n1549), .B(n1550), .Y(\iexec_stage/BUS476[2] ) );
  NAND2X2 U9 ( .A(n1556), .B(n1557), .Y(\iexec_stage/BUS476[0] ) );
  INVX2 U10 ( .A(n538), .Y(n1936) );
  AOI22XL U11 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N180 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N116 ), .B1(n855), .Y(n947) );
  CLKINVXL U12 ( .A(\iexec_stage/BUS476[4] ), .Y(n1923) );
  CLKINVXL U13 ( .A(\iexec_stage/BUS476[3] ), .Y(n574) );
  CLKINVXL U14 ( .A(\iexec_stage/BUS476[1] ), .Y(n596) );
  CLKINVXL U15 ( .A(\iexec_stage/BUS476[0] ), .Y(n597) );
  CLKINVXL U16 ( .A(\iexec_stage/BUS476[2] ), .Y(n585) );
  MXI2XL U17 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n393 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n431 ), .S0(\iexec_stage/BUS476[1] ), .Y(n109) );
  MXI2XL U18 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n391 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n429 ), .S0(\iexec_stage/BUS476[1] ), .Y(n108) );
  MXI2XL U19 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n485 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n447 ), .S0(\iexec_stage/BUS476[3] ), .Y(n103) );
  MXI2XL U20 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n485 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n515 ), .S0(\iexec_stage/BUS476[3] ), .Y(n104) );
  MXI2XL U21 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n489 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n453 ), .S0(\iexec_stage/BUS476[3] ), .Y(n105) );
  MXI2XL U22 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n489 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n519 ), .S0(\iexec_stage/BUS476[3] ), .Y(n106) );
  OAI31XL U23 ( .A0(n1927), .A1(\iexec_stage/BUS476[1] ), .A2(
        \iexec_stage/BUS476[0] ), .B0(n1926), .Y(n1469) );
  MXI2XL U24 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n368 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n372 ), .S0(\iexec_stage/BUS476[3] ), .Y(n123) );
  MXI2XL U25 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n376 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n380 ), .S0(\iexec_stage/BUS476[3] ), .Y(n124) );
  MXI2XL U26 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n557 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n545 ), .S0(\iexec_stage/BUS476[1] ), .Y(n107) );
  MXI2XL U27 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n553 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n550 ), .S0(\iexec_stage/BUS476[1] ), .Y(n112) );
  MXI2XL U28 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n586 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n590 ), .S0(\iexec_stage/BUS476[0] ), .Y(n121) );
  MXI2XL U29 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n574 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n578 ), .S0(\iexec_stage/BUS476[0] ), .Y(n118) );
  MXI2XL U30 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n578 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n582 ), .S0(\iexec_stage/BUS476[0] ), .Y(n119) );
  MXI2XL U31 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n565 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n570 ), .S0(\iexec_stage/BUS476[0] ), .Y(n113) );
  MXI2XL U32 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n562 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n546 ), .S0(\iexec_stage/BUS476[0] ), .Y(n114) );
  MXI2XL U33 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n546 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n539 ), .S0(\iexec_stage/BUS476[0] ), .Y(n115) );
  MXI2XL U34 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n539 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n565 ), .S0(\iexec_stage/BUS476[0] ), .Y(n116) );
  MXI2XL U35 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n570 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n574 ), .S0(\iexec_stage/BUS476[0] ), .Y(n117) );
  MXI2XL U36 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n582 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n586 ), .S0(\iexec_stage/BUS476[0] ), .Y(n120) );
  MXI2XL U37 ( .A(n83), .B(\iexec_stage/MIPS_alu/mips_shifter/n534 ), .S0(
        \iexec_stage/BUS476[3] ), .Y(\iexec_stage/MIPS_alu/mips_shifter/n407 )
         );
  MXI2XL U38 ( .A(\iexec_stage/BUS468[31] ), .B(\iexec_stage/BUS468[15] ), 
        .S0(\iexec_stage/BUS476[4] ), .Y(n83) );
  NAND2XL U39 ( .A(n1933), .B(n1936), .Y(n740) );
  OAI2BB2XL U40 ( .B0(n566), .B1(n565), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N112 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_0 ) );
  OAI2BB2XL U41 ( .B0(n547), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N141 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_29 ) );
  OAI2BB2XL U42 ( .B0(n543), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N116 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_4 ) );
  OAI2BB2XL U43 ( .B0(n563), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N123 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_11 ) );
  OAI2BB2XL U44 ( .B0(n542), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N117 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_5 ) );
  OAI2BB2XL U45 ( .B0(n562), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N124 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_12 ) );
  OAI2BB2XL U46 ( .B0(n541), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N118 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_6 ) );
  OAI2BB2XL U47 ( .B0(n561), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N125 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_13 ) );
  OAI2BB2XL U48 ( .B0(n540), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N119 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_7 ) );
  OAI2BB2XL U49 ( .B0(n560), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N126 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_14 ) );
  OAI2BB2XL U50 ( .B0(n539), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N120 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_8 ) );
  OAI2BB2XL U51 ( .B0(\iexec_stage/BUS468[15] ), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N127 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_15 ) );
  OAI2BB2XL U52 ( .B0(\iexec_stage/BUS468[9] ), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N121 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_9 ) );
  OAI2BB2XL U53 ( .B0(n548), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N140 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_28 ) );
  OAI2BB2XL U54 ( .B0(n549), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N139 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_27 ) );
  OAI2BB2XL U55 ( .B0(n550), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N138 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_26 ) );
  OAI2BB2XL U56 ( .B0(n551), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N137 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_25 ) );
  OAI2BB2XL U57 ( .B0(n552), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N136 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_24 ) );
  OAI2BB2XL U58 ( .B0(n553), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N135 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_23 ) );
  OAI2BB2XL U59 ( .B0(n554), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N134 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_22 ) );
  OAI2BB2XL U60 ( .B0(n555), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N133 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_21 ) );
  OAI2BB2XL U61 ( .B0(n556), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N132 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_20 ) );
  OAI2BB2XL U62 ( .B0(n557), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N131 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_19 ) );
  OAI2BB2XL U63 ( .B0(n558), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N130 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_18 ) );
  OAI2BB2XL U64 ( .B0(n559), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N129 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_17 ) );
  OAI2BB2XL U65 ( .B0(n567), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N128 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_16 ) );
  OAI2BB2XL U66 ( .B0(n564), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N122 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_10 ) );
  OAI2BB2XL U67 ( .B0(n544), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N115 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_3 ) );
  OAI2BB2XL U68 ( .B0(n546), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N114 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_2 ) );
  OAI2BB2XL U69 ( .B0(\iexec_stage/BUS468[1] ), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N113 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_1 ) );
  NAND2XL U70 ( .A(n1925), .B(\iexec_stage/BUS476[2] ), .Y(n1002) );
  OAI2BB1XL U71 ( .A0N(n565), .A1N(n597), .B0(\iexec_stage/BUS476[1] ), .Y(
        n1470) );
  OR3XL U72 ( .A(n1222), .B(\iexec_stage/BUS476[4] ), .C(n1225), .Y(n1190) );
  MXI2XL U73 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n429 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n430 ), .S0(\iexec_stage/BUS476[1] ), .Y(n110) );
  MXI2XL U74 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n481 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n530 ), .S0(\iexec_stage/BUS476[4] ), .Y(n94) );
  MXI2XL U75 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n447 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n442 ), .S0(\iexec_stage/BUS476[3] ), .Y(n96) );
  MXI2XL U76 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n468 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n465 ), .S0(\iexec_stage/BUS476[3] ), .Y(n100) );
  MXI2XL U77 ( .A(n125), .B(n126), .S0(\iexec_stage/BUS476[2] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/N195 ) );
  MXI2XL U78 ( .A(n1900), .B(n82), .S0(\iexec_stage/BUS476[0] ), .Y(n125) );
  MXI2XL U79 ( .A(n127), .B(n128), .S0(\iexec_stage/BUS476[2] ), .Y(
        \iexec_stage/MIPS_alu/mips_shifter/N194 ) );
  MXI2XL U80 ( .A(n82), .B(n1905), .S0(\iexec_stage/BUS476[0] ), .Y(n127) );
  MXI2XL U81 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n463 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n524 ), .S0(\iexec_stage/BUS476[4] ), .Y(n89) );
  MXI2XL U82 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n440 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n512 ), .S0(\iexec_stage/BUS476[4] ), .Y(n88) );
  MXI2XL U83 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n597 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n598 ), .S0(\iexec_stage/BUS476[0] ), .Y(n122) );
  MXI2XL U84 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n468 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n526 ), .S0(\iexec_stage/BUS476[3] ), .Y(n99) );
  MXI2XL U85 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n473 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n528 ), .S0(\iexec_stage/BUS476[3] ), .Y(n101) );
  MXI2XL U86 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n515 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n516 ), .S0(\iexec_stage/BUS476[3] ), .Y(n95) );
  MXI2XL U87 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n519 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n520 ), .S0(\iexec_stage/BUS476[3] ), .Y(n97) );
  OAI2BB2XL U88 ( .B0(n545), .B1(n566), .A0N(n78), .A1N(
        \iexec_stage/MIPS_alu/mips_alu/N142 ), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_30 ) );
  MXI2XL U89 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n458 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n455 ), .S0(\iexec_stage/BUS476[4] ), .Y(n91) );
  MXI2XL U90 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n493 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n383 ), .S0(\iexec_stage/BUS476[4] ), .Y(n84) );
  MXI2XL U91 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n458 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n522 ), .S0(\iexec_stage/BUS476[4] ), .Y(n92) );
  AOI22XL U92 ( .A0(cop_addr_o[24]), .A1(n1386), .B0(n1387), .B1(BUS15471[24]), 
        .Y(n1412) );
  AOI22XL U93 ( .A0(cop_addr_o[22]), .A1(n1386), .B0(n1387), .B1(BUS15471[22]), 
        .Y(n1522) );
  AOI22XL U94 ( .A0(cop_addr_o[2]), .A1(n1386), .B0(n1387), .B1(BUS15471[2]), 
        .Y(n1476) );
  AOI22XL U95 ( .A0(cop_addr_o[8]), .A1(n1386), .B0(n1387), .B1(BUS15471[8]), 
        .Y(n1487) );
  AOI22XL U96 ( .A0(cop_addr_o[21]), .A1(n1386), .B0(n1387), .B1(BUS15471[21]), 
        .Y(n1419) );
  AOI22XL U97 ( .A0(cop_addr_o[7]), .A1(n1386), .B0(n1387), .B1(BUS15471[7]), 
        .Y(n1462) );
  AOI22XL U98 ( .A0(cop_addr_o[3]), .A1(n1386), .B0(n1387), .B1(BUS15471[3]), 
        .Y(n1472) );
  AOI22XL U99 ( .A0(cop_addr_o[31]), .A1(n1386), .B0(n1387), .B1(BUS15471[31]), 
        .Y(n1540) );
  AOI22XL U100 ( .A0(cop_addr_o[11]), .A1(n1386), .B0(n1387), .B1(BUS15471[11]), .Y(n1497) );
  AOI22XL U101 ( .A0(cop_addr_o[10]), .A1(n1386), .B0(n1387), .B1(BUS15471[10]), .Y(n1492) );
  AOI22XL U102 ( .A0(cop_addr_o[20]), .A1(n1386), .B0(n1387), .B1(BUS15471[20]), .Y(n1517) );
  AOI22XL U103 ( .A0(cop_addr_o[12]), .A1(n1386), .B0(n1387), .B1(BUS15471[12]), .Y(n1450) );
  AOI22XL U104 ( .A0(cop_addr_o[19]), .A1(n1386), .B0(n1387), .B1(BUS15471[19]), .Y(n1425) );
  AOI22XL U105 ( .A0(cop_addr_o[18]), .A1(n1386), .B0(n1387), .B1(BUS15471[18]), .Y(n1431) );
  AOI22XL U106 ( .A0(cop_addr_o[13]), .A1(n1386), .B0(n1387), .B1(BUS15471[13]), .Y(n1444) );
  AOI22XL U107 ( .A0(cop_addr_o[17]), .A1(n1386), .B0(n1387), .B1(BUS15471[17]), .Y(n1512) );
  AOI22XL U108 ( .A0(cop_addr_o[15]), .A1(n1386), .B0(n1387), .B1(BUS15471[15]), .Y(n1438) );
  AOI22XL U109 ( .A0(cop_addr_o[14]), .A1(n1386), .B0(n1387), .B1(BUS15471[14]), .Y(n1502) );
  AOI22XL U110 ( .A0(cop_addr_o[16]), .A1(n1386), .B0(n1387), .B1(BUS15471[16]), .Y(n1507) );
  MXI2XL U111 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n585 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n593 ), .S0(\iexec_stage/BUS476[1] ), .Y(n82) );
  MXI2XL U112 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n560 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n557 ), .S0(\iexec_stage/BUS476[1] ), .Y(n111) );
  MXI2XL U113 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n497 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n362 ), .S0(\iexec_stage/BUS476[4] ), .Y(n85) );
  MXI2XL U114 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n501 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n468 ), .S0(\iexec_stage/BUS476[3] ), .Y(n86) );
  MXI2XL U115 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n505 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n473 ), .S0(\iexec_stage/BUS476[3] ), .Y(n87) );
  MXI2X1 U116 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n463 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n460 ), .S0(\iexec_stage/BUS476[4] ), .Y(n90) );
  MXI2X1 U117 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n481 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n478 ), .S0(\iexec_stage/BUS476[4] ), .Y(n93) );
  MXI2X1 U118 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n453 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n449 ), .S0(\iexec_stage/BUS476[3] ), .Y(n98) );
  MXI2X1 U119 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n473 ), .B(
        \iexec_stage/MIPS_alu/mips_shifter/n470 ), .S0(\iexec_stage/BUS476[3] ), .Y(n102) );
  NAND2X1 U120 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n422 ), .B(n1923), .Y(
        n126) );
  NAND2X1 U121 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n425 ), .B(n1923), .Y(
        n128) );
  INVX2 U122 ( .A(n198), .Y(n196) );
  INVX2 U123 ( .A(n198), .Y(n195) );
  INVX2 U124 ( .A(n199), .Y(n194) );
  INVX2 U125 ( .A(n199), .Y(n193) );
  INVX2 U126 ( .A(n199), .Y(n192) );
  INVX2 U127 ( .A(n200), .Y(n191) );
  INVX2 U128 ( .A(n198), .Y(n190) );
  INVX2 U129 ( .A(n199), .Y(n189) );
  INVX2 U130 ( .A(n200), .Y(n188) );
  INVX2 U131 ( .A(n198), .Y(n187) );
  INVX2 U132 ( .A(n199), .Y(n186) );
  INVX2 U133 ( .A(n199), .Y(n185) );
  INVX2 U134 ( .A(n334), .Y(n184) );
  INVX2 U135 ( .A(n334), .Y(n183) );
  INVX2 U136 ( .A(n334), .Y(n182) );
  INVX2 U137 ( .A(n200), .Y(n181) );
  INVX2 U138 ( .A(n198), .Y(n180) );
  INVX2 U139 ( .A(n200), .Y(n179) );
  INVX2 U140 ( .A(n334), .Y(n178) );
  INVX2 U141 ( .A(n200), .Y(n177) );
  INVX2 U142 ( .A(n248), .Y(n246) );
  INVX2 U143 ( .A(n248), .Y(n245) );
  INVX2 U144 ( .A(n249), .Y(n244) );
  INVX2 U145 ( .A(n249), .Y(n243) );
  INVX2 U146 ( .A(n249), .Y(n242) );
  INVX2 U147 ( .A(n250), .Y(n241) );
  INVX2 U148 ( .A(n248), .Y(n240) );
  INVX2 U149 ( .A(n249), .Y(n239) );
  INVX2 U150 ( .A(n250), .Y(n238) );
  INVX2 U151 ( .A(n248), .Y(n237) );
  INVX2 U152 ( .A(n249), .Y(n236) );
  INVX2 U153 ( .A(n249), .Y(n235) );
  INVX2 U154 ( .A(n339), .Y(n234) );
  INVX2 U155 ( .A(n339), .Y(n233) );
  INVX2 U156 ( .A(n339), .Y(n232) );
  INVX2 U157 ( .A(n250), .Y(n231) );
  INVX2 U158 ( .A(n248), .Y(n230) );
  INVX2 U159 ( .A(n250), .Y(n229) );
  INVX2 U160 ( .A(n339), .Y(n228) );
  INVX2 U161 ( .A(n250), .Y(n227) );
  INVX2 U162 ( .A(n335), .Y(n221) );
  INVX2 U163 ( .A(n335), .Y(n220) );
  INVX2 U164 ( .A(n222), .Y(n219) );
  INVX2 U165 ( .A(n222), .Y(n218) );
  INVX2 U166 ( .A(n222), .Y(n217) );
  INVX2 U167 ( .A(n223), .Y(n216) );
  INVX2 U168 ( .A(n223), .Y(n215) );
  INVX2 U169 ( .A(n223), .Y(n214) );
  INVX2 U170 ( .A(n224), .Y(n213) );
  INVX2 U171 ( .A(n224), .Y(n212) );
  INVX2 U172 ( .A(n224), .Y(n211) );
  INVX2 U173 ( .A(n225), .Y(n210) );
  INVX2 U174 ( .A(n225), .Y(n209) );
  INVX2 U175 ( .A(n225), .Y(n208) );
  INVX2 U176 ( .A(n335), .Y(n207) );
  INVX2 U177 ( .A(n222), .Y(n206) );
  INVX2 U178 ( .A(n223), .Y(n205) );
  INVX2 U179 ( .A(n223), .Y(n204) );
  INVX2 U180 ( .A(n224), .Y(n203) );
  INVX2 U181 ( .A(n225), .Y(n202) );
  INVX2 U182 ( .A(n340), .Y(n271) );
  INVX2 U183 ( .A(n340), .Y(n270) );
  INVX2 U184 ( .A(n272), .Y(n269) );
  INVX2 U185 ( .A(n272), .Y(n268) );
  INVX2 U186 ( .A(n272), .Y(n267) );
  INVX2 U187 ( .A(n273), .Y(n266) );
  INVX2 U188 ( .A(n273), .Y(n265) );
  INVX2 U189 ( .A(n273), .Y(n264) );
  INVX2 U190 ( .A(n274), .Y(n263) );
  INVX2 U191 ( .A(n274), .Y(n262) );
  INVX2 U192 ( .A(n274), .Y(n261) );
  INVX2 U193 ( .A(n275), .Y(n260) );
  INVX2 U194 ( .A(n275), .Y(n259) );
  INVX2 U195 ( .A(n275), .Y(n258) );
  INVX2 U196 ( .A(n340), .Y(n257) );
  INVX2 U197 ( .A(n272), .Y(n256) );
  INVX2 U198 ( .A(n273), .Y(n255) );
  INVX2 U199 ( .A(n273), .Y(n254) );
  INVX2 U200 ( .A(n274), .Y(n253) );
  INVX2 U201 ( .A(n275), .Y(n252) );
  INVX2 U202 ( .A(n198), .Y(n197) );
  INVX2 U203 ( .A(n248), .Y(n247) );
  INVX2 U204 ( .A(n200), .Y(n176) );
  INVX2 U205 ( .A(\iRF_stage/reg_bank/N12 ), .Y(n200) );
  INVX2 U206 ( .A(n250), .Y(n226) );
  INVX2 U207 ( .A(\iRF_stage/reg_bank/N17 ), .Y(n250) );
  INVX2 U208 ( .A(n222), .Y(n201) );
  INVX2 U209 ( .A(n272), .Y(n251) );
  INVX2 U210 ( .A(\iRF_stage/reg_bank/N12 ), .Y(n198) );
  INVX2 U211 ( .A(\iRF_stage/reg_bank/N12 ), .Y(n199) );
  INVX2 U212 ( .A(\iRF_stage/reg_bank/N13 ), .Y(n222) );
  INVX2 U213 ( .A(\iRF_stage/reg_bank/N13 ), .Y(n223) );
  INVX2 U214 ( .A(\iRF_stage/reg_bank/N13 ), .Y(n224) );
  INVX2 U215 ( .A(\iRF_stage/reg_bank/N13 ), .Y(n225) );
  INVX2 U216 ( .A(\iRF_stage/reg_bank/N17 ), .Y(n248) );
  INVX2 U217 ( .A(\iRF_stage/reg_bank/N17 ), .Y(n249) );
  INVX2 U218 ( .A(\iRF_stage/reg_bank/N18 ), .Y(n272) );
  INVX2 U219 ( .A(\iRF_stage/reg_bank/N18 ), .Y(n273) );
  INVX2 U220 ( .A(\iRF_stage/reg_bank/N18 ), .Y(n274) );
  INVX2 U221 ( .A(\iRF_stage/reg_bank/N18 ), .Y(n275) );
  OAI31X1 U222 ( .A0(n375), .A1(addr_o[1]), .A2(addr_o[0]), .B0(n376), .Y(
        wr_en_o[3]) );
  OAI21X1 U223 ( .A0(addr_o[1]), .A1(n377), .B0(n376), .Y(wr_en_o[2]) );
  OAI31X1 U224 ( .A0(n375), .A1(addr_o[0]), .A2(n378), .B0(n376), .Y(
        wr_en_o[1]) );
  NOR2X1 U225 ( .A(n379), .B(n380), .Y(n375) );
  OAI21X1 U226 ( .A0(n378), .A1(n377), .B0(n376), .Y(wr_en_o[0]) );
  NAND2X1 U227 ( .A(n379), .B(n283), .Y(n376) );
  MXI2X1 U228 ( .A(n379), .B(n380), .S0(addr_o[0]), .Y(n377) );
  CLKINVX1 U229 ( .A(n381), .Y(n380) );
  NAND3BX1 U230 ( .AN(n282), .B(n283), .C(n285), .Y(n381) );
  NOR3BX1 U231 ( .AN(n285), .B(n282), .C(n284), .Y(n379) );
  CLKINVX1 U232 ( .A(addr_o[1]), .Y(n378) );
  NAND2X1 U233 ( .A(n382), .B(n383), .Y(pc_o[9]) );
  AOI222XL U234 ( .A0(\iRF_stage/i_pc_gen/br_addr[9] ), .A1(n384), .B0(n385), 
        .B1(n54), .C0(n386), .C1(BUS7219[9]), .Y(n383) );
  AOI222XL U235 ( .A0(\iRF_stage/i_pc_gen/N43 ), .A1(n387), .B0(BUS27031[9]), 
        .B1(n388), .C0(n389), .C1(BUS24839[9]), .Y(n382) );
  NAND2X1 U236 ( .A(n390), .B(n391), .Y(pc_o[8]) );
  AOI222XL U237 ( .A0(\iRF_stage/i_pc_gen/br_addr[8] ), .A1(n384), .B0(n385), 
        .B1(n58), .C0(n386), .C1(BUS7219[8]), .Y(n391) );
  AOI222XL U238 ( .A0(\iRF_stage/i_pc_gen/N42 ), .A1(n387), .B0(BUS27031[8]), 
        .B1(n388), .C0(n389), .C1(BUS24839[8]), .Y(n390) );
  NAND2X1 U239 ( .A(n392), .B(n393), .Y(pc_o[7]) );
  AOI222XL U240 ( .A0(\iRF_stage/i_pc_gen/br_addr[7] ), .A1(n384), .B0(n385), 
        .B1(n55), .C0(n386), .C1(BUS7219[7]), .Y(n393) );
  AOI222XL U241 ( .A0(\iRF_stage/i_pc_gen/N41 ), .A1(n387), .B0(BUS27031[7]), 
        .B1(n388), .C0(n389), .C1(BUS24839[7]), .Y(n392) );
  NAND2X1 U242 ( .A(n394), .B(n395), .Y(pc_o[6]) );
  AOI222XL U243 ( .A0(\iRF_stage/i_pc_gen/br_addr[6] ), .A1(n384), .B0(n385), 
        .B1(n56), .C0(n386), .C1(BUS7219[6]), .Y(n395) );
  AOI222XL U244 ( .A0(\iRF_stage/i_pc_gen/N40 ), .A1(n387), .B0(BUS27031[6]), 
        .B1(n388), .C0(n389), .C1(BUS24839[6]), .Y(n394) );
  NAND2X1 U245 ( .A(n396), .B(n397), .Y(pc_o[5]) );
  AOI222XL U246 ( .A0(\iRF_stage/i_pc_gen/br_addr[5] ), .A1(n384), .B0(n385), 
        .B1(n57), .C0(n386), .C1(BUS7219[5]), .Y(n397) );
  AOI222XL U247 ( .A0(\iRF_stage/i_pc_gen/N39 ), .A1(n387), .B0(BUS27031[5]), 
        .B1(n388), .C0(n389), .C1(BUS24839[5]), .Y(n396) );
  NAND2X1 U248 ( .A(n398), .B(n399), .Y(pc_o[4]) );
  AOI222XL U249 ( .A0(\iRF_stage/i_pc_gen/br_addr[4] ), .A1(n384), .B0(n385), 
        .B1(n70), .C0(n386), .C1(BUS7219[4]), .Y(n399) );
  AOI222XL U250 ( .A0(\iRF_stage/i_pc_gen/N38 ), .A1(n387), .B0(BUS27031[4]), 
        .B1(n388), .C0(n389), .C1(BUS24839[4]), .Y(n398) );
  NAND2X1 U251 ( .A(n400), .B(n401), .Y(pc_o[3]) );
  AOI222XL U252 ( .A0(\iRF_stage/i_pc_gen/br_addr[3] ), .A1(n384), .B0(n385), 
        .B1(n68), .C0(n386), .C1(BUS7219[3]), .Y(n401) );
  AOI222XL U253 ( .A0(\iRF_stage/i_pc_gen/N37 ), .A1(n387), .B0(BUS27031[3]), 
        .B1(n388), .C0(n389), .C1(BUS24839[3]), .Y(n400) );
  NAND2X1 U254 ( .A(n402), .B(n403), .Y(pc_o[31]) );
  AOI222XL U255 ( .A0(\iRF_stage/i_pc_gen/br_addr[31] ), .A1(n384), .B0(
        BUS27031[31]), .B1(n404), .C0(n385), .C1(n74), .Y(n403) );
  AOI22X1 U256 ( .A0(n389), .A1(BUS24839[31]), .B0(\iRF_stage/i_pc_gen/N65 ), 
        .B1(n387), .Y(n402) );
  NAND2X1 U257 ( .A(n405), .B(n406), .Y(pc_o[30]) );
  AOI222XL U258 ( .A0(\iRF_stage/i_pc_gen/br_addr[30] ), .A1(n384), .B0(
        BUS27031[30]), .B1(n404), .C0(n385), .C1(n71), .Y(n406) );
  AOI22X1 U259 ( .A0(n389), .A1(BUS24839[30]), .B0(\iRF_stage/i_pc_gen/N64 ), 
        .B1(n387), .Y(n405) );
  OAI211X1 U260 ( .A0(n407), .A1(n408), .B0(n409), .C0(n410), .Y(pc_o[2]) );
  AOI222XL U261 ( .A0(\iRF_stage/i_pc_gen/br_addr[2] ), .A1(n384), .B0(n385), 
        .B1(n69), .C0(n386), .C1(BUS7219[2]), .Y(n410) );
  MXI2X1 U262 ( .A(n387), .B(n388), .S0(BUS27031[2]), .Y(n409) );
  NAND2X1 U263 ( .A(n411), .B(n412), .Y(pc_o[29]) );
  AOI222XL U264 ( .A0(\iRF_stage/i_pc_gen/br_addr[29] ), .A1(n384), .B0(
        BUS27031[29]), .B1(n404), .C0(n385), .C1(n72), .Y(n412) );
  AOI22X1 U265 ( .A0(n389), .A1(BUS24839[29]), .B0(\iRF_stage/i_pc_gen/N63 ), 
        .B1(n387), .Y(n411) );
  NAND2X1 U266 ( .A(n413), .B(n414), .Y(pc_o[28]) );
  AOI222XL U267 ( .A0(\iRF_stage/i_pc_gen/br_addr[28] ), .A1(n384), .B0(
        BUS27031[28]), .B1(n404), .C0(n385), .C1(n73), .Y(n414) );
  OR2X1 U268 ( .A(n388), .B(n386), .Y(n404) );
  AOI22X1 U269 ( .A0(n389), .A1(BUS24839[28]), .B0(\iRF_stage/i_pc_gen/N62 ), 
        .B1(n387), .Y(n413) );
  NAND2X1 U270 ( .A(n415), .B(n416), .Y(pc_o[27]) );
  AOI222XL U271 ( .A0(\iRF_stage/i_pc_gen/br_addr[27] ), .A1(n384), .B0(n385), 
        .B1(n45), .C0(n386), .C1(BUS7219[27]), .Y(n416) );
  AOI222XL U272 ( .A0(\iRF_stage/i_pc_gen/N61 ), .A1(n387), .B0(BUS27031[27]), 
        .B1(n388), .C0(n389), .C1(BUS24839[27]), .Y(n415) );
  NAND2X1 U273 ( .A(n417), .B(n418), .Y(pc_o[26]) );
  AOI222XL U274 ( .A0(\iRF_stage/i_pc_gen/br_addr[26] ), .A1(n384), .B0(n385), 
        .B1(n67), .C0(n386), .C1(BUS7219[26]), .Y(n418) );
  AOI222XL U275 ( .A0(\iRF_stage/i_pc_gen/N60 ), .A1(n387), .B0(BUS27031[26]), 
        .B1(n388), .C0(n389), .C1(BUS24839[26]), .Y(n417) );
  NAND2X1 U276 ( .A(n419), .B(n420), .Y(pc_o[25]) );
  AOI222XL U277 ( .A0(\iRF_stage/i_pc_gen/br_addr[25] ), .A1(n384), .B0(n385), 
        .B1(n46), .C0(n386), .C1(BUS7219[25]), .Y(n420) );
  AOI222XL U278 ( .A0(\iRF_stage/i_pc_gen/N59 ), .A1(n387), .B0(BUS27031[25]), 
        .B1(n388), .C0(n389), .C1(BUS24839[25]), .Y(n419) );
  NAND2X1 U279 ( .A(n421), .B(n422), .Y(pc_o[24]) );
  AOI222XL U280 ( .A0(\iRF_stage/i_pc_gen/br_addr[24] ), .A1(n384), .B0(n385), 
        .B1(n47), .C0(n386), .C1(BUS7219[24]), .Y(n422) );
  AOI222XL U281 ( .A0(\iRF_stage/i_pc_gen/N58 ), .A1(n387), .B0(BUS27031[24]), 
        .B1(n388), .C0(n389), .C1(BUS24839[24]), .Y(n421) );
  NAND2X1 U282 ( .A(n423), .B(n424), .Y(pc_o[23]) );
  AOI222XL U283 ( .A0(\iRF_stage/i_pc_gen/br_addr[23] ), .A1(n384), .B0(n385), 
        .B1(n66), .C0(n386), .C1(BUS7219[23]), .Y(n424) );
  AOI222XL U284 ( .A0(\iRF_stage/i_pc_gen/N57 ), .A1(n387), .B0(BUS27031[23]), 
        .B1(n388), .C0(n389), .C1(BUS24839[23]), .Y(n423) );
  NAND2X1 U285 ( .A(n425), .B(n426), .Y(pc_o[22]) );
  AOI222XL U286 ( .A0(\iRF_stage/i_pc_gen/br_addr[22] ), .A1(n384), .B0(n385), 
        .B1(n65), .C0(n386), .C1(BUS7219[22]), .Y(n426) );
  AOI222XL U287 ( .A0(\iRF_stage/i_pc_gen/N56 ), .A1(n387), .B0(BUS27031[22]), 
        .B1(n388), .C0(n389), .C1(BUS24839[22]), .Y(n425) );
  NAND2X1 U288 ( .A(n427), .B(n428), .Y(pc_o[21]) );
  AOI222XL U289 ( .A0(\iRF_stage/i_pc_gen/br_addr[21] ), .A1(n384), .B0(n385), 
        .B1(n48), .C0(n386), .C1(BUS7219[21]), .Y(n428) );
  AOI222XL U290 ( .A0(\iRF_stage/i_pc_gen/N55 ), .A1(n387), .B0(BUS27031[21]), 
        .B1(n388), .C0(n389), .C1(BUS24839[21]), .Y(n427) );
  NAND2X1 U291 ( .A(n429), .B(n430), .Y(pc_o[20]) );
  AOI222XL U292 ( .A0(\iRF_stage/i_pc_gen/br_addr[20] ), .A1(n384), .B0(n385), 
        .B1(n64), .C0(n386), .C1(BUS7219[20]), .Y(n430) );
  AOI222XL U293 ( .A0(\iRF_stage/i_pc_gen/N54 ), .A1(n387), .B0(BUS27031[20]), 
        .B1(n388), .C0(n389), .C1(BUS24839[20]), .Y(n429) );
  NAND2X1 U294 ( .A(n431), .B(n432), .Y(pc_o[1]) );
  AOI222XL U295 ( .A0(n386), .A1(BUS7219[1]), .B0(BUS27031[1]), .B1(n433), 
        .C0(n385), .C1(n75), .Y(n432) );
  AOI22X1 U296 ( .A0(\iRF_stage/i_pc_gen/br_addr[1] ), .A1(n384), .B0(n389), 
        .B1(BUS24839[1]), .Y(n431) );
  NAND2X1 U297 ( .A(n434), .B(n435), .Y(pc_o[19]) );
  AOI222XL U298 ( .A0(\iRF_stage/i_pc_gen/br_addr[19] ), .A1(n384), .B0(n385), 
        .B1(n49), .C0(n386), .C1(BUS7219[19]), .Y(n435) );
  AOI222XL U299 ( .A0(\iRF_stage/i_pc_gen/N53 ), .A1(n387), .B0(BUS27031[19]), 
        .B1(n388), .C0(n389), .C1(BUS24839[19]), .Y(n434) );
  NAND2X1 U300 ( .A(n436), .B(n437), .Y(pc_o[18]) );
  AOI222XL U301 ( .A0(\iRF_stage/i_pc_gen/br_addr[18] ), .A1(n384), .B0(n385), 
        .B1(n50), .C0(n386), .C1(BUS7219[18]), .Y(n437) );
  AOI222XL U302 ( .A0(\iRF_stage/i_pc_gen/N52 ), .A1(n387), .B0(BUS27031[18]), 
        .B1(n388), .C0(n389), .C1(BUS24839[18]), .Y(n436) );
  NAND2X1 U303 ( .A(n438), .B(n439), .Y(pc_o[17]) );
  AOI222XL U304 ( .A0(\iRF_stage/i_pc_gen/br_addr[17] ), .A1(n384), .B0(n385), 
        .B1(n63), .C0(n386), .C1(BUS7219[17]), .Y(n439) );
  AOI222XL U305 ( .A0(\iRF_stage/i_pc_gen/N51 ), .A1(n387), .B0(BUS27031[17]), 
        .B1(n388), .C0(n389), .C1(BUS24839[17]), .Y(n438) );
  NAND2X1 U306 ( .A(n440), .B(n441), .Y(pc_o[16]) );
  AOI222XL U307 ( .A0(\iRF_stage/i_pc_gen/br_addr[16] ), .A1(n384), .B0(n385), 
        .B1(n62), .C0(n386), .C1(BUS7219[16]), .Y(n441) );
  AOI222XL U308 ( .A0(\iRF_stage/i_pc_gen/N50 ), .A1(n387), .B0(BUS27031[16]), 
        .B1(n388), .C0(n389), .C1(BUS24839[16]), .Y(n440) );
  NAND2X1 U309 ( .A(n442), .B(n443), .Y(pc_o[15]) );
  AOI222XL U310 ( .A0(\iRF_stage/i_pc_gen/br_addr[15] ), .A1(n384), .B0(n385), 
        .B1(n51), .C0(n386), .C1(BUS7219[15]), .Y(n443) );
  AOI222XL U311 ( .A0(\iRF_stage/i_pc_gen/N49 ), .A1(n387), .B0(BUS27031[15]), 
        .B1(n388), .C0(n389), .C1(BUS24839[15]), .Y(n442) );
  NAND2X1 U312 ( .A(n444), .B(n445), .Y(pc_o[14]) );
  AOI222XL U313 ( .A0(\iRF_stage/i_pc_gen/br_addr[14] ), .A1(n384), .B0(n385), 
        .B1(n61), .C0(n386), .C1(BUS7219[14]), .Y(n445) );
  AOI222XL U314 ( .A0(\iRF_stage/i_pc_gen/N48 ), .A1(n387), .B0(BUS27031[14]), 
        .B1(n388), .C0(n389), .C1(BUS24839[14]), .Y(n444) );
  NAND2X1 U315 ( .A(n446), .B(n447), .Y(pc_o[13]) );
  AOI222XL U316 ( .A0(\iRF_stage/i_pc_gen/br_addr[13] ), .A1(n384), .B0(n385), 
        .B1(n52), .C0(n386), .C1(BUS7219[13]), .Y(n447) );
  AOI222XL U317 ( .A0(\iRF_stage/i_pc_gen/N47 ), .A1(n387), .B0(BUS27031[13]), 
        .B1(n388), .C0(n389), .C1(BUS24839[13]), .Y(n446) );
  NAND2X1 U318 ( .A(n448), .B(n449), .Y(pc_o[12]) );
  AOI222XL U319 ( .A0(\iRF_stage/i_pc_gen/br_addr[12] ), .A1(n384), .B0(n385), 
        .B1(n53), .C0(n386), .C1(BUS7219[12]), .Y(n449) );
  AOI222XL U320 ( .A0(\iRF_stage/i_pc_gen/N46 ), .A1(n387), .B0(BUS27031[12]), 
        .B1(n388), .C0(n389), .C1(BUS24839[12]), .Y(n448) );
  NAND2X1 U321 ( .A(n450), .B(n451), .Y(pc_o[11]) );
  AOI222XL U322 ( .A0(\iRF_stage/i_pc_gen/br_addr[11] ), .A1(n384), .B0(n385), 
        .B1(n60), .C0(n386), .C1(BUS7219[11]), .Y(n451) );
  AOI222XL U323 ( .A0(\iRF_stage/i_pc_gen/N45 ), .A1(n387), .B0(BUS27031[11]), 
        .B1(n388), .C0(n389), .C1(BUS24839[11]), .Y(n450) );
  NAND2X1 U324 ( .A(n452), .B(n453), .Y(pc_o[10]) );
  AOI222XL U325 ( .A0(\iRF_stage/i_pc_gen/br_addr[10] ), .A1(n384), .B0(n385), 
        .B1(n59), .C0(n386), .C1(BUS7219[10]), .Y(n453) );
  AOI222XL U326 ( .A0(\iRF_stage/i_pc_gen/N44 ), .A1(n387), .B0(BUS27031[10]), 
        .B1(n388), .C0(n389), .C1(BUS24839[10]), .Y(n452) );
  NAND2X1 U327 ( .A(n454), .B(n455), .Y(pc_o[0]) );
  AOI222XL U328 ( .A0(n386), .A1(BUS7219[0]), .B0(\iRF_stage/i_pc_gen/N34 ), 
        .B1(n433), .C0(n385), .C1(n76), .Y(n455) );
  NOR3BX1 U329 ( .AN(n456), .B(n302), .C(n457), .Y(n385) );
  OR2X1 U330 ( .A(n387), .B(n388), .Y(n433) );
  NOR2BX1 U331 ( .AN(n458), .B(n459), .Y(n388) );
  OAI32X1 U332 ( .A0(n460), .A1(n456), .A2(n457), .B0(n461), .B1(n462), .Y(
        n387) );
  CLKINVX1 U333 ( .A(n463), .Y(n457) );
  OR2X1 U334 ( .A(n464), .B(n465), .Y(n460) );
  AND2X1 U335 ( .A(n465), .B(n463), .Y(n386) );
  AND3X2 U336 ( .A(n302), .B(n38), .C(n303), .Y(n465) );
  AOI22X1 U337 ( .A0(\iRF_stage/i_pc_gen/br_addr[0] ), .A1(n384), .B0(n389), 
        .B1(BUS24839[0]), .Y(n454) );
  CLKINVX1 U338 ( .A(n408), .Y(n389) );
  NAND2X1 U339 ( .A(n464), .B(n463), .Y(n408) );
  NOR3BX1 U340 ( .AN(n303), .B(n38), .C(n302), .Y(n464) );
  NOR2BX1 U341 ( .AN(n462), .B(n461), .Y(n384) );
  NAND3X1 U342 ( .A(n463), .B(n456), .C(n302), .Y(n461) );
  NOR2X1 U343 ( .A(n38), .B(n303), .Y(n456) );
  AOI2BB1X1 U344 ( .A0N(n1935), .A1N(n466), .B0(n467), .Y(n463) );
  MX2X1 U345 ( .A(n468), .B(n469), .S0(n295), .Y(n462) );
  OAI2BB1X1 U346 ( .A0N(n470), .A1N(n293), .B0(n471), .Y(n469) );
  MXI2X1 U347 ( .A(n472), .B(n473), .S0(n294), .Y(n471) );
  CLKINVX1 U348 ( .A(n470), .Y(n473) );
  NOR2X1 U349 ( .A(n293), .B(n474), .Y(n472) );
  NAND2X1 U350 ( .A(n475), .B(n476), .Y(n470) );
  NOR4X1 U351 ( .A(n477), .B(n478), .C(n479), .D(n480), .Y(n476) );
  NAND4X1 U352 ( .A(n481), .B(n482), .C(n483), .D(n484), .Y(n480) );
  XNOR2X1 U353 ( .A(BUS7160[20]), .B(BUS24839[20]), .Y(n484) );
  XNOR2X1 U354 ( .A(BUS7160[21]), .B(BUS24839[21]), .Y(n483) );
  XNOR2X1 U355 ( .A(BUS7160[22]), .B(BUS24839[22]), .Y(n482) );
  XNOR2X1 U356 ( .A(BUS7160[23]), .B(BUS24839[23]), .Y(n481) );
  NAND4X1 U357 ( .A(n485), .B(n486), .C(n487), .D(n488), .Y(n479) );
  XNOR2X1 U358 ( .A(BUS7160[17]), .B(BUS24839[17]), .Y(n488) );
  XNOR2X1 U359 ( .A(BUS7160[18]), .B(BUS24839[18]), .Y(n487) );
  XNOR2X1 U360 ( .A(BUS7160[19]), .B(BUS24839[19]), .Y(n486) );
  XNOR2X1 U361 ( .A(BUS7160[1]), .B(BUS24839[1]), .Y(n485) );
  NAND4X1 U362 ( .A(n489), .B(n490), .C(n491), .D(n492), .Y(n478) );
  XNOR2X1 U363 ( .A(BUS7160[13]), .B(BUS24839[13]), .Y(n492) );
  XNOR2X1 U364 ( .A(BUS7160[14]), .B(BUS24839[14]), .Y(n491) );
  XNOR2X1 U365 ( .A(BUS7160[15]), .B(BUS24839[15]), .Y(n490) );
  XNOR2X1 U366 ( .A(BUS7160[16]), .B(BUS24839[16]), .Y(n489) );
  NAND4X1 U367 ( .A(n493), .B(n494), .C(n495), .D(n496), .Y(n477) );
  XOR2X1 U368 ( .A(BUS7160[0]), .B(n497), .Y(n496) );
  XOR2X1 U369 ( .A(BUS7160[10]), .B(n498), .Y(n495) );
  XOR2X1 U370 ( .A(BUS7160[11]), .B(n499), .Y(n494) );
  XNOR2X1 U371 ( .A(BUS7160[12]), .B(BUS24839[12]), .Y(n493) );
  NOR4X1 U372 ( .A(n500), .B(n501), .C(n502), .D(n503), .Y(n475) );
  NAND4X1 U373 ( .A(n504), .B(n505), .C(n506), .D(n507), .Y(n503) );
  XNOR2X1 U374 ( .A(BUS7160[6]), .B(BUS24839[6]), .Y(n507) );
  XNOR2X1 U375 ( .A(BUS7160[7]), .B(BUS24839[7]), .Y(n506) );
  XNOR2X1 U376 ( .A(BUS7160[8]), .B(BUS24839[8]), .Y(n505) );
  XNOR2X1 U377 ( .A(BUS7160[9]), .B(BUS24839[9]), .Y(n504) );
  NAND4X1 U378 ( .A(n508), .B(n509), .C(n510), .D(n511), .Y(n502) );
  XOR2X1 U379 ( .A(BUS7160[31]), .B(n512), .Y(n511) );
  XNOR2X1 U380 ( .A(BUS7160[3]), .B(BUS24839[3]), .Y(n510) );
  XNOR2X1 U381 ( .A(BUS7160[4]), .B(BUS24839[4]), .Y(n509) );
  XNOR2X1 U382 ( .A(BUS7160[5]), .B(BUS24839[5]), .Y(n508) );
  NAND4X1 U383 ( .A(n513), .B(n514), .C(n515), .D(n516), .Y(n501) );
  XNOR2X1 U384 ( .A(BUS7160[28]), .B(BUS24839[28]), .Y(n516) );
  XNOR2X1 U385 ( .A(BUS7160[29]), .B(BUS24839[29]), .Y(n515) );
  XOR2X1 U386 ( .A(BUS7160[2]), .B(n407), .Y(n514) );
  CLKINVX1 U387 ( .A(BUS24839[2]), .Y(n407) );
  XNOR2X1 U388 ( .A(BUS7160[30]), .B(BUS24839[30]), .Y(n513) );
  NAND4X1 U389 ( .A(n517), .B(n518), .C(n519), .D(n520), .Y(n500) );
  XNOR2X1 U390 ( .A(BUS7160[24]), .B(BUS24839[24]), .Y(n520) );
  XNOR2X1 U391 ( .A(BUS7160[25]), .B(BUS24839[25]), .Y(n519) );
  XNOR2X1 U392 ( .A(BUS7160[26]), .B(BUS24839[26]), .Y(n518) );
  XNOR2X1 U393 ( .A(BUS7160[27]), .B(BUS24839[27]), .Y(n517) );
  OAI21X1 U394 ( .A0(n294), .A1(n512), .B0(n521), .Y(n468) );
  MXI2X1 U395 ( .A(n474), .B(n522), .S0(n293), .Y(n521) );
  AND2X1 U396 ( .A(n512), .B(n294), .Y(n522) );
  CLKINVX1 U397 ( .A(n523), .Y(n474) );
  OAI31X1 U398 ( .A0(n524), .A1(n525), .A2(n526), .B0(n512), .Y(n523) );
  NAND4X1 U399 ( .A(n498), .B(n499), .C(n497), .D(n527), .Y(n526) );
  NOR4X1 U400 ( .A(BUS24839[15]), .B(BUS24839[14]), .C(BUS24839[13]), .D(
        BUS24839[12]), .Y(n527) );
  CLKINVX1 U401 ( .A(BUS24839[0]), .Y(n497) );
  CLKINVX1 U402 ( .A(BUS24839[11]), .Y(n499) );
  CLKINVX1 U403 ( .A(BUS24839[10]), .Y(n498) );
  NAND2X1 U404 ( .A(n528), .B(n529), .Y(n525) );
  NOR4X1 U405 ( .A(BUS24839[22]), .B(BUS24839[21]), .C(BUS24839[20]), .D(
        BUS24839[1]), .Y(n529) );
  NOR4X1 U406 ( .A(BUS24839[19]), .B(BUS24839[18]), .C(BUS24839[17]), .D(
        BUS24839[16]), .Y(n528) );
  NAND4X1 U407 ( .A(n530), .B(n531), .C(n532), .D(n533), .Y(n524) );
  NOR4X1 U408 ( .A(BUS24839[9]), .B(BUS24839[8]), .C(BUS24839[7]), .D(
        BUS24839[6]), .Y(n533) );
  NOR4X1 U409 ( .A(BUS24839[5]), .B(BUS24839[4]), .C(BUS24839[3]), .D(
        BUS24839[30]), .Y(n532) );
  NOR4X1 U410 ( .A(BUS24839[2]), .B(BUS24839[29]), .C(BUS24839[28]), .D(
        BUS24839[27]), .Y(n531) );
  NOR4X1 U411 ( .A(BUS24839[26]), .B(BUS24839[25]), .C(BUS24839[24]), .D(
        BUS24839[23]), .Y(n530) );
  CLKINVX1 U412 ( .A(BUS24839[31]), .Y(n512) );
  CLKINVX1 U413 ( .A(addr_o[31]), .Y(n1878) );
  OAI2BB1X1 U414 ( .A0N(n78), .A1N(\iexec_stage/MIPS_alu/mips_alu/N143 ), .B0(
        n534), .Y(n1879) );
  CLKINVX1 U415 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n477 ), .Y(n1880) );
  CLKINVX1 U416 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n362 ), .Y(n1882) );
  CLKINVX1 U417 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n553 ), .Y(n1884) );
  CLKINVX1 U418 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n383 ), .Y(n1887) );
  CLKINVX1 U419 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n562 ), .Y(n1888) );
  CLKINVX1 U420 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n440 ), .Y(n1890) );
  CLKINVX1 U421 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n386 ), .Y(n1894) );
  CLKINVX1 U422 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n590 ), .Y(n1900) );
  CLKINVX1 U423 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n585 ), .Y(n1902) );
  CLKINVX1 U424 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n589 ), .Y(n1904) );
  CLKINVX1 U425 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n597 ), .Y(n1905) );
  CLKINVX1 U426 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n390 ), .Y(n1907) );
  CLKINVX1 U427 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n392 ), .Y(n1908) );
  CLKINVX1 U428 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n391 ), .Y(n1910) );
  CLKINVX1 U429 ( .A(\iexec_stage/MIPS_alu/mips_shifter/n431 ), .Y(n1914) );
  OAI21X1 U430 ( .A0(n535), .A1(n536), .B0(n1936), .Y(n1929) );
  CLKINVX1 U431 ( .A(n537), .Y(n1930) );
  NOR2X1 U432 ( .A(iack_o), .B(n538), .Y(n1932) );
  NOR2X1 U433 ( .A(n538), .B(n467), .Y(n1934) );
  CLKINVX1 U434 ( .A(BUS27031[2]), .Y(n1939) );
  XOR2X1 U435 ( .A(\iexec_stage/BUS468[9] ), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[9] ) );
  XOR2X1 U436 ( .A(n539), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[8] ) );
  XOR2X1 U437 ( .A(n540), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[7] ) );
  XOR2X1 U438 ( .A(n541), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[6] ) );
  XOR2X1 U439 ( .A(n542), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[5] ) );
  XOR2X1 U440 ( .A(n543), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[4] ) );
  XOR2X1 U441 ( .A(n544), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[3] ) );
  XOR2X1 U442 ( .A(\iexec_stage/BUS468[31] ), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[31] ) );
  XOR2X1 U443 ( .A(n545), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[30] ) );
  XOR2X1 U444 ( .A(n546), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[2] ) );
  XOR2X1 U445 ( .A(n547), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[29] ) );
  XOR2X1 U446 ( .A(n548), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[28] ) );
  XOR2X1 U447 ( .A(n549), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[27] ) );
  XOR2X1 U448 ( .A(n550), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[26] ) );
  XOR2X1 U449 ( .A(n551), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[25] ) );
  XOR2X1 U450 ( .A(n552), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[24] ) );
  XOR2X1 U451 ( .A(n553), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[23] ) );
  XOR2X1 U452 ( .A(n554), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[22] ) );
  XOR2X1 U453 ( .A(n555), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[21] ) );
  XOR2X1 U454 ( .A(n556), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[20] ) );
  XOR2X1 U455 ( .A(\iexec_stage/BUS468[1] ), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[1] ) );
  XOR2X1 U456 ( .A(n557), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[19] ) );
  XOR2X1 U457 ( .A(n558), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[18] ) );
  XOR2X1 U458 ( .A(n559), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[17] ) );
  XOR2X1 U459 ( .A(n1), .B(n1906), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[16] ) );
  XOR2X1 U460 ( .A(\iexec_stage/BUS468[15] ), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[15] ) );
  XOR2X1 U461 ( .A(n560), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[14] ) );
  XOR2X1 U462 ( .A(n561), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[13] ) );
  XOR2X1 U463 ( .A(n562), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[12] ) );
  XOR2X1 U464 ( .A(n563), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[11] ) );
  XOR2X1 U465 ( .A(n564), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[10] ) );
  XOR2X1 U466 ( .A(n565), .B(n78), .Y(
        \iexec_stage/MIPS_alu/mips_alu/r92/B_AS[0] ) );
  CLKINVX1 U467 ( .A(n534), .Y(\iexec_stage/MIPS_alu/mips_alu/U3/U3/Z_32 ) );
  NAND2X1 U468 ( .A(n1938), .B(n1881), .Y(n534) );
  NOR2X1 U469 ( .A(n568), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_9 ) );
  NOR2X1 U470 ( .A(n569), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_8 ) );
  NOR2X1 U471 ( .A(n570), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_7 ) );
  NOR2X1 U472 ( .A(n571), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_6 ) );
  NOR2X1 U473 ( .A(n572), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_5 ) );
  NOR2X1 U474 ( .A(n1923), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_4 ) );
  NOR2X1 U475 ( .A(n573), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_32 ) );
  AND2X1 U476 ( .A(\iexec_stage/BUS476[30] ), .B(n1938), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_30 ) );
  NOR2X1 U477 ( .A(n574), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_3 ) );
  NOR2X1 U478 ( .A(n575), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_29 ) );
  NOR2X1 U479 ( .A(n576), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_28 ) );
  NOR2X1 U480 ( .A(n577), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_27 ) );
  NOR2X1 U481 ( .A(n578), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_26 ) );
  NOR2X1 U482 ( .A(n579), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_25 ) );
  NOR2X1 U483 ( .A(n580), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_24 ) );
  NOR2X1 U484 ( .A(n581), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_23 ) );
  NOR2X1 U485 ( .A(n582), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_22 ) );
  NOR2X1 U486 ( .A(n583), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_21 ) );
  NOR2X1 U487 ( .A(n584), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_20 ) );
  NOR2X1 U488 ( .A(n585), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_2 ) );
  NOR2X1 U489 ( .A(n586), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_19 ) );
  NOR2X1 U490 ( .A(n587), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_18 ) );
  NOR2X1 U491 ( .A(n588), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_17 ) );
  NOR2X1 U492 ( .A(n589), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_16 ) );
  NOR2X1 U493 ( .A(n590), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_15 ) );
  NOR2X1 U494 ( .A(n591), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_14 ) );
  NOR2X1 U495 ( .A(n592), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_13 ) );
  NOR2X1 U496 ( .A(n593), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_12 ) );
  NOR2X1 U497 ( .A(n594), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_11 ) );
  NOR2X1 U498 ( .A(n595), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_10 ) );
  NOR2X1 U499 ( .A(n596), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_1 ) );
  NOR2X1 U500 ( .A(n597), .B(n566), .Y(
        \iexec_stage/MIPS_alu/mips_alu/U3/U2/Z_0 ) );
  CLKINVX1 U501 ( .A(n1938), .Y(n566) );
  OAI21X1 U502 ( .A0(n1935), .A1(n304), .B0(n598), .Y(iack_o) );
  MX2X1 U503 ( .A(\iRF_stage/reg_bank/reg_bank[861] ), .B(n13), .S0(n599), .Y(
        \iRF_stage/reg_bank/n999 ) );
  MX2X1 U504 ( .A(\iRF_stage/reg_bank/reg_bank[860] ), .B(n14), .S0(n599), .Y(
        \iRF_stage/reg_bank/n998 ) );
  MX2X1 U505 ( .A(\iRF_stage/reg_bank/reg_bank[859] ), .B(n15), .S0(n599), .Y(
        \iRF_stage/reg_bank/n997 ) );
  MX2X1 U506 ( .A(\iRF_stage/reg_bank/reg_bank[858] ), .B(n16), .S0(n599), .Y(
        \iRF_stage/reg_bank/n996 ) );
  MX2X1 U507 ( .A(\iRF_stage/reg_bank/reg_bank[857] ), .B(n17), .S0(n599), .Y(
        \iRF_stage/reg_bank/n995 ) );
  MX2X1 U508 ( .A(\iRF_stage/reg_bank/reg_bank[856] ), .B(n18), .S0(n599), .Y(
        \iRF_stage/reg_bank/n994 ) );
  MX2X1 U509 ( .A(\iRF_stage/reg_bank/reg_bank[855] ), .B(n19), .S0(n599), .Y(
        \iRF_stage/reg_bank/n993 ) );
  MX2X1 U510 ( .A(\iRF_stage/reg_bank/reg_bank[854] ), .B(n20), .S0(n599), .Y(
        \iRF_stage/reg_bank/n992 ) );
  MX2X1 U511 ( .A(\iRF_stage/reg_bank/reg_bank[853] ), .B(n21), .S0(n599), .Y(
        \iRF_stage/reg_bank/n991 ) );
  MX2X1 U512 ( .A(\iRF_stage/reg_bank/reg_bank[852] ), .B(n22), .S0(n599), .Y(
        \iRF_stage/reg_bank/n990 ) );
  MX2X1 U513 ( .A(\iRF_stage/reg_bank/reg_bank[851] ), .B(n24), .S0(n599), .Y(
        \iRF_stage/reg_bank/n989 ) );
  MX2X1 U514 ( .A(\iRF_stage/reg_bank/reg_bank[850] ), .B(n25), .S0(n599), .Y(
        \iRF_stage/reg_bank/n988 ) );
  MX2X1 U515 ( .A(\iRF_stage/reg_bank/reg_bank[849] ), .B(n26), .S0(n599), .Y(
        \iRF_stage/reg_bank/n987 ) );
  MX2X1 U516 ( .A(\iRF_stage/reg_bank/reg_bank[848] ), .B(n27), .S0(n599), .Y(
        \iRF_stage/reg_bank/n986 ) );
  MX2X1 U517 ( .A(\iRF_stage/reg_bank/reg_bank[847] ), .B(n28), .S0(n599), .Y(
        \iRF_stage/reg_bank/n985 ) );
  MX2X1 U518 ( .A(\iRF_stage/reg_bank/reg_bank[846] ), .B(n29), .S0(n599), .Y(
        \iRF_stage/reg_bank/n984 ) );
  MX2X1 U519 ( .A(\iRF_stage/reg_bank/reg_bank[845] ), .B(n30), .S0(n599), .Y(
        \iRF_stage/reg_bank/n983 ) );
  MX2X1 U520 ( .A(\iRF_stage/reg_bank/reg_bank[844] ), .B(n31), .S0(n599), .Y(
        \iRF_stage/reg_bank/n982 ) );
  MX2X1 U521 ( .A(\iRF_stage/reg_bank/reg_bank[843] ), .B(n32), .S0(n599), .Y(
        \iRF_stage/reg_bank/n981 ) );
  MX2X1 U522 ( .A(\iRF_stage/reg_bank/reg_bank[842] ), .B(n33), .S0(n599), .Y(
        \iRF_stage/reg_bank/n980 ) );
  MX2X1 U523 ( .A(\iRF_stage/reg_bank/reg_bank[841] ), .B(n3), .S0(n599), .Y(
        \iRF_stage/reg_bank/n979 ) );
  MX2X1 U524 ( .A(\iRF_stage/reg_bank/reg_bank[840] ), .B(n4), .S0(n599), .Y(
        \iRF_stage/reg_bank/n978 ) );
  MX2X1 U525 ( .A(\iRF_stage/reg_bank/reg_bank[839] ), .B(n5), .S0(n599), .Y(
        \iRF_stage/reg_bank/n977 ) );
  MX2X1 U526 ( .A(\iRF_stage/reg_bank/reg_bank[838] ), .B(n6), .S0(n599), .Y(
        \iRF_stage/reg_bank/n976 ) );
  MX2X1 U527 ( .A(\iRF_stage/reg_bank/reg_bank[837] ), .B(n7), .S0(n599), .Y(
        \iRF_stage/reg_bank/n975 ) );
  MX2X1 U528 ( .A(\iRF_stage/reg_bank/reg_bank[836] ), .B(n8), .S0(n599), .Y(
        \iRF_stage/reg_bank/n974 ) );
  MX2X1 U529 ( .A(\iRF_stage/reg_bank/reg_bank[835] ), .B(n9), .S0(n599), .Y(
        \iRF_stage/reg_bank/n973 ) );
  MX2X1 U530 ( .A(\iRF_stage/reg_bank/reg_bank[834] ), .B(n12), .S0(n599), .Y(
        \iRF_stage/reg_bank/n972 ) );
  MX2X1 U531 ( .A(\iRF_stage/reg_bank/reg_bank[833] ), .B(n23), .S0(n599), .Y(
        \iRF_stage/reg_bank/n971 ) );
  MX2X1 U532 ( .A(\iRF_stage/reg_bank/reg_bank[832] ), .B(n34), .S0(n599), .Y(
        \iRF_stage/reg_bank/n970 ) );
  MX2X1 U533 ( .A(\iRF_stage/reg_bank/reg_bank[831] ), .B(n10), .S0(n600), .Y(
        \iRF_stage/reg_bank/n969 ) );
  MX2X1 U534 ( .A(\iRF_stage/reg_bank/reg_bank[830] ), .B(n11), .S0(n600), .Y(
        \iRF_stage/reg_bank/n968 ) );
  MX2X1 U535 ( .A(\iRF_stage/reg_bank/reg_bank[829] ), .B(n13), .S0(n600), .Y(
        \iRF_stage/reg_bank/n967 ) );
  MX2X1 U536 ( .A(\iRF_stage/reg_bank/reg_bank[828] ), .B(n14), .S0(n600), .Y(
        \iRF_stage/reg_bank/n966 ) );
  MX2X1 U537 ( .A(\iRF_stage/reg_bank/reg_bank[827] ), .B(n15), .S0(n600), .Y(
        \iRF_stage/reg_bank/n965 ) );
  MX2X1 U538 ( .A(\iRF_stage/reg_bank/reg_bank[826] ), .B(n16), .S0(n600), .Y(
        \iRF_stage/reg_bank/n964 ) );
  MX2X1 U539 ( .A(\iRF_stage/reg_bank/reg_bank[825] ), .B(n17), .S0(n600), .Y(
        \iRF_stage/reg_bank/n963 ) );
  MX2X1 U540 ( .A(\iRF_stage/reg_bank/reg_bank[824] ), .B(n18), .S0(n600), .Y(
        \iRF_stage/reg_bank/n962 ) );
  MX2X1 U541 ( .A(\iRF_stage/reg_bank/reg_bank[823] ), .B(n19), .S0(n600), .Y(
        \iRF_stage/reg_bank/n961 ) );
  MX2X1 U542 ( .A(\iRF_stage/reg_bank/reg_bank[822] ), .B(n20), .S0(n600), .Y(
        \iRF_stage/reg_bank/n960 ) );
  MX2X1 U543 ( .A(\iRF_stage/reg_bank/reg_bank[821] ), .B(n21), .S0(n600), .Y(
        \iRF_stage/reg_bank/n959 ) );
  MX2X1 U544 ( .A(\iRF_stage/reg_bank/reg_bank[820] ), .B(n22), .S0(n600), .Y(
        \iRF_stage/reg_bank/n958 ) );
  MX2X1 U545 ( .A(\iRF_stage/reg_bank/reg_bank[819] ), .B(n24), .S0(n600), .Y(
        \iRF_stage/reg_bank/n957 ) );
  MX2X1 U546 ( .A(\iRF_stage/reg_bank/reg_bank[818] ), .B(n25), .S0(n600), .Y(
        \iRF_stage/reg_bank/n956 ) );
  MX2X1 U547 ( .A(\iRF_stage/reg_bank/reg_bank[817] ), .B(n26), .S0(n600), .Y(
        \iRF_stage/reg_bank/n955 ) );
  MX2X1 U548 ( .A(\iRF_stage/reg_bank/reg_bank[816] ), .B(n27), .S0(n600), .Y(
        \iRF_stage/reg_bank/n954 ) );
  MX2X1 U549 ( .A(\iRF_stage/reg_bank/reg_bank[815] ), .B(n28), .S0(n600), .Y(
        \iRF_stage/reg_bank/n953 ) );
  MX2X1 U550 ( .A(\iRF_stage/reg_bank/reg_bank[814] ), .B(n29), .S0(n600), .Y(
        \iRF_stage/reg_bank/n952 ) );
  MX2X1 U551 ( .A(\iRF_stage/reg_bank/reg_bank[813] ), .B(n30), .S0(n600), .Y(
        \iRF_stage/reg_bank/n951 ) );
  MX2X1 U552 ( .A(\iRF_stage/reg_bank/reg_bank[812] ), .B(n31), .S0(n600), .Y(
        \iRF_stage/reg_bank/n950 ) );
  MX2X1 U553 ( .A(\iRF_stage/reg_bank/reg_bank[811] ), .B(n32), .S0(n600), .Y(
        \iRF_stage/reg_bank/n949 ) );
  MX2X1 U554 ( .A(\iRF_stage/reg_bank/reg_bank[810] ), .B(n33), .S0(n600), .Y(
        \iRF_stage/reg_bank/n948 ) );
  MX2X1 U555 ( .A(\iRF_stage/reg_bank/reg_bank[809] ), .B(n3), .S0(n600), .Y(
        \iRF_stage/reg_bank/n947 ) );
  MX2X1 U556 ( .A(\iRF_stage/reg_bank/reg_bank[808] ), .B(n4), .S0(n600), .Y(
        \iRF_stage/reg_bank/n946 ) );
  MX2X1 U557 ( .A(\iRF_stage/reg_bank/reg_bank[807] ), .B(n5), .S0(n600), .Y(
        \iRF_stage/reg_bank/n945 ) );
  MX2X1 U558 ( .A(\iRF_stage/reg_bank/reg_bank[806] ), .B(n6), .S0(n600), .Y(
        \iRF_stage/reg_bank/n944 ) );
  MX2X1 U559 ( .A(\iRF_stage/reg_bank/reg_bank[805] ), .B(n7), .S0(n600), .Y(
        \iRF_stage/reg_bank/n943 ) );
  MX2X1 U560 ( .A(\iRF_stage/reg_bank/reg_bank[804] ), .B(n8), .S0(n600), .Y(
        \iRF_stage/reg_bank/n942 ) );
  MX2X1 U561 ( .A(\iRF_stage/reg_bank/reg_bank[803] ), .B(n9), .S0(n600), .Y(
        \iRF_stage/reg_bank/n941 ) );
  MX2X1 U562 ( .A(\iRF_stage/reg_bank/reg_bank[802] ), .B(n12), .S0(n600), .Y(
        \iRF_stage/reg_bank/n940 ) );
  MX2X1 U563 ( .A(\iRF_stage/reg_bank/reg_bank[801] ), .B(n23), .S0(n600), .Y(
        \iRF_stage/reg_bank/n939 ) );
  MX2X1 U564 ( .A(\iRF_stage/reg_bank/reg_bank[800] ), .B(n34), .S0(n600), .Y(
        \iRF_stage/reg_bank/n938 ) );
  AND2X1 U565 ( .A(n601), .B(n602), .Y(n600) );
  MX2X1 U566 ( .A(\iRF_stage/reg_bank/reg_bank[799] ), .B(n10), .S0(n603), .Y(
        \iRF_stage/reg_bank/n937 ) );
  MX2X1 U567 ( .A(\iRF_stage/reg_bank/reg_bank[798] ), .B(n11), .S0(n603), .Y(
        \iRF_stage/reg_bank/n936 ) );
  MX2X1 U568 ( .A(\iRF_stage/reg_bank/reg_bank[797] ), .B(n13), .S0(n603), .Y(
        \iRF_stage/reg_bank/n935 ) );
  MX2X1 U569 ( .A(\iRF_stage/reg_bank/reg_bank[796] ), .B(n14), .S0(n603), .Y(
        \iRF_stage/reg_bank/n934 ) );
  MX2X1 U570 ( .A(\iRF_stage/reg_bank/reg_bank[795] ), .B(n15), .S0(n603), .Y(
        \iRF_stage/reg_bank/n933 ) );
  MX2X1 U571 ( .A(\iRF_stage/reg_bank/reg_bank[794] ), .B(n16), .S0(n603), .Y(
        \iRF_stage/reg_bank/n932 ) );
  MX2X1 U572 ( .A(\iRF_stage/reg_bank/reg_bank[793] ), .B(n17), .S0(n603), .Y(
        \iRF_stage/reg_bank/n931 ) );
  MX2X1 U573 ( .A(\iRF_stage/reg_bank/reg_bank[792] ), .B(n18), .S0(n603), .Y(
        \iRF_stage/reg_bank/n930 ) );
  MX2X1 U574 ( .A(\iRF_stage/reg_bank/reg_bank[791] ), .B(n19), .S0(n603), .Y(
        \iRF_stage/reg_bank/n929 ) );
  MX2X1 U575 ( .A(\iRF_stage/reg_bank/reg_bank[790] ), .B(n20), .S0(n603), .Y(
        \iRF_stage/reg_bank/n928 ) );
  MX2X1 U576 ( .A(\iRF_stage/reg_bank/reg_bank[789] ), .B(n21), .S0(n603), .Y(
        \iRF_stage/reg_bank/n927 ) );
  MX2X1 U577 ( .A(\iRF_stage/reg_bank/reg_bank[788] ), .B(n22), .S0(n603), .Y(
        \iRF_stage/reg_bank/n926 ) );
  MX2X1 U578 ( .A(\iRF_stage/reg_bank/reg_bank[787] ), .B(n24), .S0(n603), .Y(
        \iRF_stage/reg_bank/n925 ) );
  MX2X1 U579 ( .A(\iRF_stage/reg_bank/reg_bank[786] ), .B(n25), .S0(n603), .Y(
        \iRF_stage/reg_bank/n924 ) );
  MX2X1 U580 ( .A(\iRF_stage/reg_bank/reg_bank[785] ), .B(n26), .S0(n603), .Y(
        \iRF_stage/reg_bank/n923 ) );
  MX2X1 U581 ( .A(\iRF_stage/reg_bank/reg_bank[784] ), .B(n27), .S0(n603), .Y(
        \iRF_stage/reg_bank/n922 ) );
  MX2X1 U582 ( .A(\iRF_stage/reg_bank/reg_bank[783] ), .B(n28), .S0(n603), .Y(
        \iRF_stage/reg_bank/n921 ) );
  MX2X1 U583 ( .A(\iRF_stage/reg_bank/reg_bank[782] ), .B(n29), .S0(n603), .Y(
        \iRF_stage/reg_bank/n920 ) );
  MX2X1 U584 ( .A(\iRF_stage/reg_bank/reg_bank[781] ), .B(n30), .S0(n603), .Y(
        \iRF_stage/reg_bank/n919 ) );
  MX2X1 U585 ( .A(\iRF_stage/reg_bank/reg_bank[780] ), .B(n31), .S0(n603), .Y(
        \iRF_stage/reg_bank/n918 ) );
  MX2X1 U586 ( .A(\iRF_stage/reg_bank/reg_bank[779] ), .B(n32), .S0(n603), .Y(
        \iRF_stage/reg_bank/n917 ) );
  MX2X1 U587 ( .A(\iRF_stage/reg_bank/reg_bank[778] ), .B(n33), .S0(n603), .Y(
        \iRF_stage/reg_bank/n916 ) );
  MX2X1 U588 ( .A(\iRF_stage/reg_bank/reg_bank[777] ), .B(n3), .S0(n603), .Y(
        \iRF_stage/reg_bank/n915 ) );
  MX2X1 U589 ( .A(\iRF_stage/reg_bank/reg_bank[776] ), .B(n4), .S0(n603), .Y(
        \iRF_stage/reg_bank/n914 ) );
  MX2X1 U590 ( .A(\iRF_stage/reg_bank/reg_bank[775] ), .B(n5), .S0(n603), .Y(
        \iRF_stage/reg_bank/n913 ) );
  MX2X1 U591 ( .A(\iRF_stage/reg_bank/reg_bank[774] ), .B(n6), .S0(n603), .Y(
        \iRF_stage/reg_bank/n912 ) );
  MX2X1 U592 ( .A(\iRF_stage/reg_bank/reg_bank[773] ), .B(n7), .S0(n603), .Y(
        \iRF_stage/reg_bank/n911 ) );
  MX2X1 U593 ( .A(\iRF_stage/reg_bank/reg_bank[772] ), .B(n8), .S0(n603), .Y(
        \iRF_stage/reg_bank/n910 ) );
  MX2X1 U594 ( .A(\iRF_stage/reg_bank/reg_bank[771] ), .B(n9), .S0(n603), .Y(
        \iRF_stage/reg_bank/n909 ) );
  MX2X1 U595 ( .A(\iRF_stage/reg_bank/reg_bank[770] ), .B(n12), .S0(n603), .Y(
        \iRF_stage/reg_bank/n908 ) );
  MX2X1 U596 ( .A(\iRF_stage/reg_bank/reg_bank[769] ), .B(n23), .S0(n603), .Y(
        \iRF_stage/reg_bank/n907 ) );
  MX2X1 U597 ( .A(\iRF_stage/reg_bank/reg_bank[768] ), .B(n34), .S0(n603), .Y(
        \iRF_stage/reg_bank/n906 ) );
  AND2X1 U598 ( .A(n604), .B(n602), .Y(n603) );
  MX2X1 U599 ( .A(\iRF_stage/reg_bank/reg_bank[767] ), .B(n10), .S0(n605), .Y(
        \iRF_stage/reg_bank/n905 ) );
  MX2X1 U600 ( .A(\iRF_stage/reg_bank/reg_bank[766] ), .B(n11), .S0(n605), .Y(
        \iRF_stage/reg_bank/n904 ) );
  MX2X1 U601 ( .A(\iRF_stage/reg_bank/reg_bank[765] ), .B(n13), .S0(n605), .Y(
        \iRF_stage/reg_bank/n903 ) );
  MX2X1 U602 ( .A(\iRF_stage/reg_bank/reg_bank[764] ), .B(n14), .S0(n605), .Y(
        \iRF_stage/reg_bank/n902 ) );
  MX2X1 U603 ( .A(\iRF_stage/reg_bank/reg_bank[763] ), .B(n15), .S0(n605), .Y(
        \iRF_stage/reg_bank/n901 ) );
  MX2X1 U604 ( .A(\iRF_stage/reg_bank/reg_bank[762] ), .B(n16), .S0(n605), .Y(
        \iRF_stage/reg_bank/n900 ) );
  MX2X1 U605 ( .A(\iRF_stage/reg_bank/reg_bank[761] ), .B(n17), .S0(n605), .Y(
        \iRF_stage/reg_bank/n899 ) );
  MX2X1 U606 ( .A(\iRF_stage/reg_bank/reg_bank[760] ), .B(n18), .S0(n605), .Y(
        \iRF_stage/reg_bank/n898 ) );
  MX2X1 U607 ( .A(\iRF_stage/reg_bank/reg_bank[759] ), .B(n19), .S0(n605), .Y(
        \iRF_stage/reg_bank/n897 ) );
  MX2X1 U608 ( .A(\iRF_stage/reg_bank/reg_bank[758] ), .B(n20), .S0(n605), .Y(
        \iRF_stage/reg_bank/n896 ) );
  MX2X1 U609 ( .A(\iRF_stage/reg_bank/reg_bank[757] ), .B(n21), .S0(n605), .Y(
        \iRF_stage/reg_bank/n895 ) );
  MX2X1 U610 ( .A(\iRF_stage/reg_bank/reg_bank[756] ), .B(n22), .S0(n605), .Y(
        \iRF_stage/reg_bank/n894 ) );
  MX2X1 U611 ( .A(\iRF_stage/reg_bank/reg_bank[755] ), .B(n24), .S0(n605), .Y(
        \iRF_stage/reg_bank/n893 ) );
  MX2X1 U612 ( .A(\iRF_stage/reg_bank/reg_bank[754] ), .B(n25), .S0(n605), .Y(
        \iRF_stage/reg_bank/n892 ) );
  MX2X1 U613 ( .A(\iRF_stage/reg_bank/reg_bank[753] ), .B(n26), .S0(n605), .Y(
        \iRF_stage/reg_bank/n891 ) );
  MX2X1 U614 ( .A(\iRF_stage/reg_bank/reg_bank[752] ), .B(n27), .S0(n605), .Y(
        \iRF_stage/reg_bank/n890 ) );
  MX2X1 U615 ( .A(\iRF_stage/reg_bank/reg_bank[751] ), .B(n28), .S0(n605), .Y(
        \iRF_stage/reg_bank/n889 ) );
  MX2X1 U616 ( .A(\iRF_stage/reg_bank/reg_bank[750] ), .B(n29), .S0(n605), .Y(
        \iRF_stage/reg_bank/n888 ) );
  MX2X1 U617 ( .A(\iRF_stage/reg_bank/reg_bank[749] ), .B(n30), .S0(n605), .Y(
        \iRF_stage/reg_bank/n887 ) );
  MX2X1 U618 ( .A(\iRF_stage/reg_bank/reg_bank[748] ), .B(n31), .S0(n605), .Y(
        \iRF_stage/reg_bank/n886 ) );
  MX2X1 U619 ( .A(\iRF_stage/reg_bank/reg_bank[747] ), .B(n32), .S0(n605), .Y(
        \iRF_stage/reg_bank/n885 ) );
  MX2X1 U620 ( .A(\iRF_stage/reg_bank/reg_bank[746] ), .B(n33), .S0(n605), .Y(
        \iRF_stage/reg_bank/n884 ) );
  MX2X1 U621 ( .A(\iRF_stage/reg_bank/reg_bank[745] ), .B(n3), .S0(n605), .Y(
        \iRF_stage/reg_bank/n883 ) );
  MX2X1 U622 ( .A(\iRF_stage/reg_bank/reg_bank[744] ), .B(n4), .S0(n605), .Y(
        \iRF_stage/reg_bank/n882 ) );
  MX2X1 U623 ( .A(\iRF_stage/reg_bank/reg_bank[743] ), .B(n5), .S0(n605), .Y(
        \iRF_stage/reg_bank/n881 ) );
  MX2X1 U624 ( .A(\iRF_stage/reg_bank/reg_bank[742] ), .B(n6), .S0(n605), .Y(
        \iRF_stage/reg_bank/n880 ) );
  MX2X1 U625 ( .A(\iRF_stage/reg_bank/reg_bank[741] ), .B(n7), .S0(n605), .Y(
        \iRF_stage/reg_bank/n879 ) );
  MX2X1 U626 ( .A(\iRF_stage/reg_bank/reg_bank[740] ), .B(n8), .S0(n605), .Y(
        \iRF_stage/reg_bank/n878 ) );
  MX2X1 U627 ( .A(\iRF_stage/reg_bank/reg_bank[739] ), .B(n9), .S0(n605), .Y(
        \iRF_stage/reg_bank/n877 ) );
  MX2X1 U628 ( .A(\iRF_stage/reg_bank/reg_bank[738] ), .B(n12), .S0(n605), .Y(
        \iRF_stage/reg_bank/n876 ) );
  MX2X1 U629 ( .A(\iRF_stage/reg_bank/reg_bank[737] ), .B(n23), .S0(n605), .Y(
        \iRF_stage/reg_bank/n875 ) );
  MX2X1 U630 ( .A(\iRF_stage/reg_bank/reg_bank[736] ), .B(n34), .S0(n605), .Y(
        \iRF_stage/reg_bank/n874 ) );
  AND2X1 U631 ( .A(n606), .B(n607), .Y(n605) );
  MX2X1 U632 ( .A(\iRF_stage/reg_bank/reg_bank[735] ), .B(n10), .S0(n608), .Y(
        \iRF_stage/reg_bank/n873 ) );
  MX2X1 U633 ( .A(\iRF_stage/reg_bank/reg_bank[734] ), .B(n11), .S0(n608), .Y(
        \iRF_stage/reg_bank/n872 ) );
  MX2X1 U634 ( .A(\iRF_stage/reg_bank/reg_bank[733] ), .B(n13), .S0(n608), .Y(
        \iRF_stage/reg_bank/n871 ) );
  MX2X1 U635 ( .A(\iRF_stage/reg_bank/reg_bank[732] ), .B(n14), .S0(n608), .Y(
        \iRF_stage/reg_bank/n870 ) );
  MX2X1 U636 ( .A(\iRF_stage/reg_bank/reg_bank[731] ), .B(n15), .S0(n608), .Y(
        \iRF_stage/reg_bank/n869 ) );
  MX2X1 U637 ( .A(\iRF_stage/reg_bank/reg_bank[730] ), .B(n16), .S0(n608), .Y(
        \iRF_stage/reg_bank/n868 ) );
  MX2X1 U638 ( .A(\iRF_stage/reg_bank/reg_bank[729] ), .B(n17), .S0(n608), .Y(
        \iRF_stage/reg_bank/n867 ) );
  MX2X1 U639 ( .A(\iRF_stage/reg_bank/reg_bank[728] ), .B(n18), .S0(n608), .Y(
        \iRF_stage/reg_bank/n866 ) );
  MX2X1 U640 ( .A(\iRF_stage/reg_bank/reg_bank[727] ), .B(n19), .S0(n608), .Y(
        \iRF_stage/reg_bank/n865 ) );
  MX2X1 U641 ( .A(\iRF_stage/reg_bank/reg_bank[726] ), .B(n20), .S0(n608), .Y(
        \iRF_stage/reg_bank/n864 ) );
  MX2X1 U642 ( .A(\iRF_stage/reg_bank/reg_bank[725] ), .B(n21), .S0(n608), .Y(
        \iRF_stage/reg_bank/n863 ) );
  MX2X1 U643 ( .A(\iRF_stage/reg_bank/reg_bank[724] ), .B(n22), .S0(n608), .Y(
        \iRF_stage/reg_bank/n862 ) );
  MX2X1 U644 ( .A(\iRF_stage/reg_bank/reg_bank[723] ), .B(n24), .S0(n608), .Y(
        \iRF_stage/reg_bank/n861 ) );
  MX2X1 U645 ( .A(\iRF_stage/reg_bank/reg_bank[722] ), .B(n25), .S0(n608), .Y(
        \iRF_stage/reg_bank/n860 ) );
  MX2X1 U646 ( .A(\iRF_stage/reg_bank/reg_bank[721] ), .B(n26), .S0(n608), .Y(
        \iRF_stage/reg_bank/n859 ) );
  MX2X1 U647 ( .A(\iRF_stage/reg_bank/reg_bank[720] ), .B(n27), .S0(n608), .Y(
        \iRF_stage/reg_bank/n858 ) );
  MX2X1 U648 ( .A(\iRF_stage/reg_bank/reg_bank[719] ), .B(n28), .S0(n608), .Y(
        \iRF_stage/reg_bank/n857 ) );
  MX2X1 U649 ( .A(\iRF_stage/reg_bank/reg_bank[718] ), .B(n29), .S0(n608), .Y(
        \iRF_stage/reg_bank/n856 ) );
  MX2X1 U650 ( .A(\iRF_stage/reg_bank/reg_bank[717] ), .B(n30), .S0(n608), .Y(
        \iRF_stage/reg_bank/n855 ) );
  MX2X1 U651 ( .A(\iRF_stage/reg_bank/reg_bank[716] ), .B(n31), .S0(n608), .Y(
        \iRF_stage/reg_bank/n854 ) );
  MX2X1 U652 ( .A(\iRF_stage/reg_bank/reg_bank[715] ), .B(n32), .S0(n608), .Y(
        \iRF_stage/reg_bank/n853 ) );
  MX2X1 U653 ( .A(\iRF_stage/reg_bank/reg_bank[714] ), .B(n33), .S0(n608), .Y(
        \iRF_stage/reg_bank/n852 ) );
  MX2X1 U654 ( .A(\iRF_stage/reg_bank/reg_bank[713] ), .B(n3), .S0(n608), .Y(
        \iRF_stage/reg_bank/n851 ) );
  MX2X1 U655 ( .A(\iRF_stage/reg_bank/reg_bank[712] ), .B(n4), .S0(n608), .Y(
        \iRF_stage/reg_bank/n850 ) );
  MX2X1 U656 ( .A(\iRF_stage/reg_bank/reg_bank[711] ), .B(n5), .S0(n608), .Y(
        \iRF_stage/reg_bank/n849 ) );
  MX2X1 U657 ( .A(\iRF_stage/reg_bank/reg_bank[710] ), .B(n6), .S0(n608), .Y(
        \iRF_stage/reg_bank/n848 ) );
  MX2X1 U658 ( .A(\iRF_stage/reg_bank/reg_bank[709] ), .B(n7), .S0(n608), .Y(
        \iRF_stage/reg_bank/n847 ) );
  MX2X1 U659 ( .A(\iRF_stage/reg_bank/reg_bank[708] ), .B(n8), .S0(n608), .Y(
        \iRF_stage/reg_bank/n846 ) );
  MX2X1 U660 ( .A(\iRF_stage/reg_bank/reg_bank[707] ), .B(n9), .S0(n608), .Y(
        \iRF_stage/reg_bank/n845 ) );
  MX2X1 U661 ( .A(\iRF_stage/reg_bank/reg_bank[706] ), .B(n12), .S0(n608), .Y(
        \iRF_stage/reg_bank/n844 ) );
  MX2X1 U662 ( .A(\iRF_stage/reg_bank/reg_bank[705] ), .B(n23), .S0(n608), .Y(
        \iRF_stage/reg_bank/n843 ) );
  MX2X1 U663 ( .A(\iRF_stage/reg_bank/reg_bank[704] ), .B(n34), .S0(n608), .Y(
        \iRF_stage/reg_bank/n842 ) );
  AND2X1 U664 ( .A(n609), .B(n607), .Y(n608) );
  MX2X1 U665 ( .A(\iRF_stage/reg_bank/reg_bank[703] ), .B(n10), .S0(n610), .Y(
        \iRF_stage/reg_bank/n841 ) );
  MX2X1 U666 ( .A(\iRF_stage/reg_bank/reg_bank[702] ), .B(n11), .S0(n610), .Y(
        \iRF_stage/reg_bank/n840 ) );
  MX2X1 U667 ( .A(\iRF_stage/reg_bank/reg_bank[701] ), .B(n13), .S0(n610), .Y(
        \iRF_stage/reg_bank/n839 ) );
  MX2X1 U668 ( .A(\iRF_stage/reg_bank/reg_bank[700] ), .B(n14), .S0(n610), .Y(
        \iRF_stage/reg_bank/n838 ) );
  MX2X1 U669 ( .A(\iRF_stage/reg_bank/reg_bank[699] ), .B(n15), .S0(n610), .Y(
        \iRF_stage/reg_bank/n837 ) );
  MX2X1 U670 ( .A(\iRF_stage/reg_bank/reg_bank[698] ), .B(n16), .S0(n610), .Y(
        \iRF_stage/reg_bank/n836 ) );
  MX2X1 U671 ( .A(\iRF_stage/reg_bank/reg_bank[697] ), .B(n17), .S0(n610), .Y(
        \iRF_stage/reg_bank/n835 ) );
  MX2X1 U672 ( .A(\iRF_stage/reg_bank/reg_bank[696] ), .B(n18), .S0(n610), .Y(
        \iRF_stage/reg_bank/n834 ) );
  MX2X1 U673 ( .A(\iRF_stage/reg_bank/reg_bank[695] ), .B(n19), .S0(n610), .Y(
        \iRF_stage/reg_bank/n833 ) );
  MX2X1 U674 ( .A(\iRF_stage/reg_bank/reg_bank[694] ), .B(n20), .S0(n610), .Y(
        \iRF_stage/reg_bank/n832 ) );
  MX2X1 U675 ( .A(\iRF_stage/reg_bank/reg_bank[693] ), .B(n21), .S0(n610), .Y(
        \iRF_stage/reg_bank/n831 ) );
  MX2X1 U676 ( .A(\iRF_stage/reg_bank/reg_bank[692] ), .B(n22), .S0(n610), .Y(
        \iRF_stage/reg_bank/n830 ) );
  MX2X1 U677 ( .A(\iRF_stage/reg_bank/reg_bank[691] ), .B(n24), .S0(n610), .Y(
        \iRF_stage/reg_bank/n829 ) );
  MX2X1 U678 ( .A(\iRF_stage/reg_bank/reg_bank[690] ), .B(n25), .S0(n610), .Y(
        \iRF_stage/reg_bank/n828 ) );
  MX2X1 U679 ( .A(\iRF_stage/reg_bank/reg_bank[689] ), .B(n26), .S0(n610), .Y(
        \iRF_stage/reg_bank/n827 ) );
  MX2X1 U680 ( .A(\iRF_stage/reg_bank/reg_bank[688] ), .B(n27), .S0(n610), .Y(
        \iRF_stage/reg_bank/n826 ) );
  MX2X1 U681 ( .A(\iRF_stage/reg_bank/reg_bank[687] ), .B(n28), .S0(n610), .Y(
        \iRF_stage/reg_bank/n825 ) );
  MX2X1 U682 ( .A(\iRF_stage/reg_bank/reg_bank[686] ), .B(n29), .S0(n610), .Y(
        \iRF_stage/reg_bank/n824 ) );
  MX2X1 U683 ( .A(\iRF_stage/reg_bank/reg_bank[685] ), .B(n30), .S0(n610), .Y(
        \iRF_stage/reg_bank/n823 ) );
  MX2X1 U684 ( .A(\iRF_stage/reg_bank/reg_bank[684] ), .B(n31), .S0(n610), .Y(
        \iRF_stage/reg_bank/n822 ) );
  MX2X1 U685 ( .A(\iRF_stage/reg_bank/reg_bank[683] ), .B(n32), .S0(n610), .Y(
        \iRF_stage/reg_bank/n821 ) );
  MX2X1 U686 ( .A(\iRF_stage/reg_bank/reg_bank[682] ), .B(n33), .S0(n610), .Y(
        \iRF_stage/reg_bank/n820 ) );
  MX2X1 U687 ( .A(\iRF_stage/reg_bank/reg_bank[681] ), .B(n3), .S0(n610), .Y(
        \iRF_stage/reg_bank/n819 ) );
  MX2X1 U688 ( .A(\iRF_stage/reg_bank/reg_bank[680] ), .B(n4), .S0(n610), .Y(
        \iRF_stage/reg_bank/n818 ) );
  MX2X1 U689 ( .A(\iRF_stage/reg_bank/reg_bank[679] ), .B(n5), .S0(n610), .Y(
        \iRF_stage/reg_bank/n817 ) );
  MX2X1 U690 ( .A(\iRF_stage/reg_bank/reg_bank[678] ), .B(n6), .S0(n610), .Y(
        \iRF_stage/reg_bank/n816 ) );
  MX2X1 U691 ( .A(\iRF_stage/reg_bank/reg_bank[677] ), .B(n7), .S0(n610), .Y(
        \iRF_stage/reg_bank/n815 ) );
  MX2X1 U692 ( .A(\iRF_stage/reg_bank/reg_bank[676] ), .B(n8), .S0(n610), .Y(
        \iRF_stage/reg_bank/n814 ) );
  MX2X1 U693 ( .A(\iRF_stage/reg_bank/reg_bank[675] ), .B(n9), .S0(n610), .Y(
        \iRF_stage/reg_bank/n813 ) );
  MX2X1 U694 ( .A(\iRF_stage/reg_bank/reg_bank[674] ), .B(n12), .S0(n610), .Y(
        \iRF_stage/reg_bank/n812 ) );
  MX2X1 U695 ( .A(\iRF_stage/reg_bank/reg_bank[673] ), .B(n23), .S0(n610), .Y(
        \iRF_stage/reg_bank/n811 ) );
  MX2X1 U696 ( .A(\iRF_stage/reg_bank/reg_bank[672] ), .B(n34), .S0(n610), .Y(
        \iRF_stage/reg_bank/n810 ) );
  AND2X1 U697 ( .A(n611), .B(n607), .Y(n610) );
  MX2X1 U698 ( .A(\iRF_stage/reg_bank/reg_bank[671] ), .B(n10), .S0(n612), .Y(
        \iRF_stage/reg_bank/n809 ) );
  MX2X1 U699 ( .A(\iRF_stage/reg_bank/reg_bank[670] ), .B(n11), .S0(n612), .Y(
        \iRF_stage/reg_bank/n808 ) );
  MX2X1 U700 ( .A(\iRF_stage/reg_bank/reg_bank[669] ), .B(n13), .S0(n612), .Y(
        \iRF_stage/reg_bank/n807 ) );
  MX2X1 U701 ( .A(\iRF_stage/reg_bank/reg_bank[668] ), .B(n14), .S0(n612), .Y(
        \iRF_stage/reg_bank/n806 ) );
  MX2X1 U702 ( .A(\iRF_stage/reg_bank/reg_bank[667] ), .B(n15), .S0(n612), .Y(
        \iRF_stage/reg_bank/n805 ) );
  MX2X1 U703 ( .A(\iRF_stage/reg_bank/reg_bank[666] ), .B(n16), .S0(n612), .Y(
        \iRF_stage/reg_bank/n804 ) );
  MX2X1 U704 ( .A(\iRF_stage/reg_bank/reg_bank[665] ), .B(n17), .S0(n612), .Y(
        \iRF_stage/reg_bank/n803 ) );
  MX2X1 U705 ( .A(\iRF_stage/reg_bank/reg_bank[664] ), .B(n18), .S0(n612), .Y(
        \iRF_stage/reg_bank/n802 ) );
  MX2X1 U706 ( .A(\iRF_stage/reg_bank/reg_bank[663] ), .B(n19), .S0(n612), .Y(
        \iRF_stage/reg_bank/n801 ) );
  MX2X1 U707 ( .A(\iRF_stage/reg_bank/reg_bank[662] ), .B(n20), .S0(n612), .Y(
        \iRF_stage/reg_bank/n800 ) );
  MX2X1 U708 ( .A(\iRF_stage/reg_bank/reg_bank[661] ), .B(n21), .S0(n612), .Y(
        \iRF_stage/reg_bank/n799 ) );
  MX2X1 U709 ( .A(\iRF_stage/reg_bank/reg_bank[660] ), .B(n22), .S0(n612), .Y(
        \iRF_stage/reg_bank/n798 ) );
  MX2X1 U710 ( .A(\iRF_stage/reg_bank/reg_bank[659] ), .B(n24), .S0(n612), .Y(
        \iRF_stage/reg_bank/n797 ) );
  MX2X1 U711 ( .A(\iRF_stage/reg_bank/reg_bank[658] ), .B(n25), .S0(n612), .Y(
        \iRF_stage/reg_bank/n796 ) );
  MX2X1 U712 ( .A(\iRF_stage/reg_bank/reg_bank[657] ), .B(n26), .S0(n612), .Y(
        \iRF_stage/reg_bank/n795 ) );
  MX2X1 U713 ( .A(\iRF_stage/reg_bank/reg_bank[656] ), .B(n27), .S0(n612), .Y(
        \iRF_stage/reg_bank/n794 ) );
  MX2X1 U714 ( .A(\iRF_stage/reg_bank/reg_bank[655] ), .B(n28), .S0(n612), .Y(
        \iRF_stage/reg_bank/n793 ) );
  MX2X1 U715 ( .A(\iRF_stage/reg_bank/reg_bank[654] ), .B(n29), .S0(n612), .Y(
        \iRF_stage/reg_bank/n792 ) );
  MX2X1 U716 ( .A(\iRF_stage/reg_bank/reg_bank[653] ), .B(n30), .S0(n612), .Y(
        \iRF_stage/reg_bank/n791 ) );
  MX2X1 U717 ( .A(\iRF_stage/reg_bank/reg_bank[652] ), .B(n31), .S0(n612), .Y(
        \iRF_stage/reg_bank/n790 ) );
  MX2X1 U718 ( .A(\iRF_stage/reg_bank/reg_bank[651] ), .B(n32), .S0(n612), .Y(
        \iRF_stage/reg_bank/n789 ) );
  MX2X1 U719 ( .A(\iRF_stage/reg_bank/reg_bank[650] ), .B(n33), .S0(n612), .Y(
        \iRF_stage/reg_bank/n788 ) );
  MX2X1 U720 ( .A(\iRF_stage/reg_bank/reg_bank[649] ), .B(n3), .S0(n612), .Y(
        \iRF_stage/reg_bank/n787 ) );
  MX2X1 U721 ( .A(\iRF_stage/reg_bank/reg_bank[648] ), .B(n4), .S0(n612), .Y(
        \iRF_stage/reg_bank/n786 ) );
  MX2X1 U722 ( .A(\iRF_stage/reg_bank/reg_bank[647] ), .B(n5), .S0(n612), .Y(
        \iRF_stage/reg_bank/n785 ) );
  MX2X1 U723 ( .A(\iRF_stage/reg_bank/reg_bank[646] ), .B(n6), .S0(n612), .Y(
        \iRF_stage/reg_bank/n784 ) );
  MX2X1 U724 ( .A(\iRF_stage/reg_bank/reg_bank[645] ), .B(n7), .S0(n612), .Y(
        \iRF_stage/reg_bank/n783 ) );
  MX2X1 U725 ( .A(\iRF_stage/reg_bank/reg_bank[644] ), .B(n8), .S0(n612), .Y(
        \iRF_stage/reg_bank/n782 ) );
  MX2X1 U726 ( .A(\iRF_stage/reg_bank/reg_bank[643] ), .B(n9), .S0(n612), .Y(
        \iRF_stage/reg_bank/n781 ) );
  MX2X1 U727 ( .A(\iRF_stage/reg_bank/reg_bank[642] ), .B(n12), .S0(n612), .Y(
        \iRF_stage/reg_bank/n780 ) );
  MX2X1 U728 ( .A(\iRF_stage/reg_bank/reg_bank[641] ), .B(n23), .S0(n612), .Y(
        \iRF_stage/reg_bank/n779 ) );
  MX2X1 U729 ( .A(\iRF_stage/reg_bank/reg_bank[640] ), .B(n34), .S0(n612), .Y(
        \iRF_stage/reg_bank/n778 ) );
  AND2X1 U730 ( .A(n613), .B(n607), .Y(n612) );
  MX2X1 U731 ( .A(\iRF_stage/reg_bank/reg_bank[639] ), .B(n10), .S0(n614), .Y(
        \iRF_stage/reg_bank/n777 ) );
  MX2X1 U732 ( .A(\iRF_stage/reg_bank/reg_bank[638] ), .B(n11), .S0(n614), .Y(
        \iRF_stage/reg_bank/n776 ) );
  MX2X1 U733 ( .A(\iRF_stage/reg_bank/reg_bank[637] ), .B(n13), .S0(n614), .Y(
        \iRF_stage/reg_bank/n775 ) );
  MX2X1 U734 ( .A(\iRF_stage/reg_bank/reg_bank[636] ), .B(n14), .S0(n614), .Y(
        \iRF_stage/reg_bank/n774 ) );
  MX2X1 U735 ( .A(\iRF_stage/reg_bank/reg_bank[635] ), .B(n15), .S0(n614), .Y(
        \iRF_stage/reg_bank/n773 ) );
  MX2X1 U736 ( .A(\iRF_stage/reg_bank/reg_bank[634] ), .B(n16), .S0(n614), .Y(
        \iRF_stage/reg_bank/n772 ) );
  MX2X1 U737 ( .A(\iRF_stage/reg_bank/reg_bank[633] ), .B(n17), .S0(n614), .Y(
        \iRF_stage/reg_bank/n771 ) );
  MX2X1 U738 ( .A(\iRF_stage/reg_bank/reg_bank[632] ), .B(n18), .S0(n614), .Y(
        \iRF_stage/reg_bank/n770 ) );
  MX2X1 U739 ( .A(\iRF_stage/reg_bank/reg_bank[631] ), .B(n19), .S0(n614), .Y(
        \iRF_stage/reg_bank/n769 ) );
  MX2X1 U740 ( .A(\iRF_stage/reg_bank/reg_bank[630] ), .B(n20), .S0(n614), .Y(
        \iRF_stage/reg_bank/n768 ) );
  MX2X1 U741 ( .A(\iRF_stage/reg_bank/reg_bank[629] ), .B(n21), .S0(n614), .Y(
        \iRF_stage/reg_bank/n767 ) );
  MX2X1 U742 ( .A(\iRF_stage/reg_bank/reg_bank[628] ), .B(n22), .S0(n614), .Y(
        \iRF_stage/reg_bank/n766 ) );
  MX2X1 U743 ( .A(\iRF_stage/reg_bank/reg_bank[627] ), .B(n24), .S0(n614), .Y(
        \iRF_stage/reg_bank/n765 ) );
  MX2X1 U744 ( .A(\iRF_stage/reg_bank/reg_bank[626] ), .B(n25), .S0(n614), .Y(
        \iRF_stage/reg_bank/n764 ) );
  MX2X1 U745 ( .A(\iRF_stage/reg_bank/reg_bank[625] ), .B(n26), .S0(n614), .Y(
        \iRF_stage/reg_bank/n763 ) );
  MX2X1 U746 ( .A(\iRF_stage/reg_bank/reg_bank[624] ), .B(n27), .S0(n614), .Y(
        \iRF_stage/reg_bank/n762 ) );
  MX2X1 U747 ( .A(\iRF_stage/reg_bank/reg_bank[623] ), .B(n28), .S0(n614), .Y(
        \iRF_stage/reg_bank/n761 ) );
  MX2X1 U748 ( .A(\iRF_stage/reg_bank/reg_bank[622] ), .B(n29), .S0(n614), .Y(
        \iRF_stage/reg_bank/n760 ) );
  MX2X1 U749 ( .A(\iRF_stage/reg_bank/reg_bank[621] ), .B(n30), .S0(n614), .Y(
        \iRF_stage/reg_bank/n759 ) );
  MX2X1 U750 ( .A(\iRF_stage/reg_bank/reg_bank[620] ), .B(n31), .S0(n614), .Y(
        \iRF_stage/reg_bank/n758 ) );
  MX2X1 U751 ( .A(\iRF_stage/reg_bank/reg_bank[619] ), .B(n32), .S0(n614), .Y(
        \iRF_stage/reg_bank/n757 ) );
  MX2X1 U752 ( .A(\iRF_stage/reg_bank/reg_bank[618] ), .B(n33), .S0(n614), .Y(
        \iRF_stage/reg_bank/n756 ) );
  MX2X1 U753 ( .A(\iRF_stage/reg_bank/reg_bank[617] ), .B(n3), .S0(n614), .Y(
        \iRF_stage/reg_bank/n755 ) );
  MX2X1 U754 ( .A(\iRF_stage/reg_bank/reg_bank[616] ), .B(n4), .S0(n614), .Y(
        \iRF_stage/reg_bank/n754 ) );
  MX2X1 U755 ( .A(\iRF_stage/reg_bank/reg_bank[615] ), .B(n5), .S0(n614), .Y(
        \iRF_stage/reg_bank/n753 ) );
  MX2X1 U756 ( .A(\iRF_stage/reg_bank/reg_bank[614] ), .B(n6), .S0(n614), .Y(
        \iRF_stage/reg_bank/n752 ) );
  MX2X1 U757 ( .A(\iRF_stage/reg_bank/reg_bank[613] ), .B(n7), .S0(n614), .Y(
        \iRF_stage/reg_bank/n751 ) );
  MX2X1 U758 ( .A(\iRF_stage/reg_bank/reg_bank[612] ), .B(n8), .S0(n614), .Y(
        \iRF_stage/reg_bank/n750 ) );
  MX2X1 U759 ( .A(\iRF_stage/reg_bank/reg_bank[611] ), .B(n9), .S0(n614), .Y(
        \iRF_stage/reg_bank/n749 ) );
  MX2X1 U760 ( .A(\iRF_stage/reg_bank/reg_bank[610] ), .B(n12), .S0(n614), .Y(
        \iRF_stage/reg_bank/n748 ) );
  MX2X1 U761 ( .A(\iRF_stage/reg_bank/reg_bank[609] ), .B(n23), .S0(n614), .Y(
        \iRF_stage/reg_bank/n747 ) );
  MX2X1 U762 ( .A(\iRF_stage/reg_bank/reg_bank[608] ), .B(n34), .S0(n614), .Y(
        \iRF_stage/reg_bank/n746 ) );
  AND2X1 U763 ( .A(n615), .B(n607), .Y(n614) );
  MX2X1 U764 ( .A(\iRF_stage/reg_bank/reg_bank[607] ), .B(n10), .S0(n616), .Y(
        \iRF_stage/reg_bank/n745 ) );
  MX2X1 U765 ( .A(\iRF_stage/reg_bank/reg_bank[606] ), .B(n11), .S0(n616), .Y(
        \iRF_stage/reg_bank/n744 ) );
  MX2X1 U766 ( .A(\iRF_stage/reg_bank/reg_bank[605] ), .B(n13), .S0(n616), .Y(
        \iRF_stage/reg_bank/n743 ) );
  MX2X1 U767 ( .A(\iRF_stage/reg_bank/reg_bank[604] ), .B(n14), .S0(n616), .Y(
        \iRF_stage/reg_bank/n742 ) );
  MX2X1 U768 ( .A(\iRF_stage/reg_bank/reg_bank[603] ), .B(n15), .S0(n616), .Y(
        \iRF_stage/reg_bank/n741 ) );
  MX2X1 U769 ( .A(\iRF_stage/reg_bank/reg_bank[602] ), .B(n16), .S0(n616), .Y(
        \iRF_stage/reg_bank/n740 ) );
  MX2X1 U770 ( .A(\iRF_stage/reg_bank/reg_bank[601] ), .B(n17), .S0(n616), .Y(
        \iRF_stage/reg_bank/n739 ) );
  MX2X1 U771 ( .A(\iRF_stage/reg_bank/reg_bank[600] ), .B(n18), .S0(n616), .Y(
        \iRF_stage/reg_bank/n738 ) );
  MX2X1 U772 ( .A(\iRF_stage/reg_bank/reg_bank[599] ), .B(n19), .S0(n616), .Y(
        \iRF_stage/reg_bank/n737 ) );
  MX2X1 U773 ( .A(\iRF_stage/reg_bank/reg_bank[598] ), .B(n20), .S0(n616), .Y(
        \iRF_stage/reg_bank/n736 ) );
  MX2X1 U774 ( .A(\iRF_stage/reg_bank/reg_bank[597] ), .B(n21), .S0(n616), .Y(
        \iRF_stage/reg_bank/n735 ) );
  MX2X1 U775 ( .A(\iRF_stage/reg_bank/reg_bank[596] ), .B(n22), .S0(n616), .Y(
        \iRF_stage/reg_bank/n734 ) );
  MX2X1 U776 ( .A(\iRF_stage/reg_bank/reg_bank[595] ), .B(n24), .S0(n616), .Y(
        \iRF_stage/reg_bank/n733 ) );
  MX2X1 U777 ( .A(\iRF_stage/reg_bank/reg_bank[594] ), .B(n25), .S0(n616), .Y(
        \iRF_stage/reg_bank/n732 ) );
  MX2X1 U778 ( .A(\iRF_stage/reg_bank/reg_bank[593] ), .B(n26), .S0(n616), .Y(
        \iRF_stage/reg_bank/n731 ) );
  MX2X1 U779 ( .A(\iRF_stage/reg_bank/reg_bank[592] ), .B(n27), .S0(n616), .Y(
        \iRF_stage/reg_bank/n730 ) );
  MX2X1 U780 ( .A(\iRF_stage/reg_bank/reg_bank[591] ), .B(n28), .S0(n616), .Y(
        \iRF_stage/reg_bank/n729 ) );
  MX2X1 U781 ( .A(\iRF_stage/reg_bank/reg_bank[590] ), .B(n29), .S0(n616), .Y(
        \iRF_stage/reg_bank/n728 ) );
  MX2X1 U782 ( .A(\iRF_stage/reg_bank/reg_bank[589] ), .B(n30), .S0(n616), .Y(
        \iRF_stage/reg_bank/n727 ) );
  MX2X1 U783 ( .A(\iRF_stage/reg_bank/reg_bank[588] ), .B(n31), .S0(n616), .Y(
        \iRF_stage/reg_bank/n726 ) );
  MX2X1 U784 ( .A(\iRF_stage/reg_bank/reg_bank[587] ), .B(n32), .S0(n616), .Y(
        \iRF_stage/reg_bank/n725 ) );
  MX2X1 U785 ( .A(\iRF_stage/reg_bank/reg_bank[586] ), .B(n33), .S0(n616), .Y(
        \iRF_stage/reg_bank/n724 ) );
  MX2X1 U786 ( .A(\iRF_stage/reg_bank/reg_bank[585] ), .B(n3), .S0(n616), .Y(
        \iRF_stage/reg_bank/n723 ) );
  MX2X1 U787 ( .A(\iRF_stage/reg_bank/reg_bank[584] ), .B(n4), .S0(n616), .Y(
        \iRF_stage/reg_bank/n722 ) );
  MX2X1 U788 ( .A(\iRF_stage/reg_bank/reg_bank[583] ), .B(n5), .S0(n616), .Y(
        \iRF_stage/reg_bank/n721 ) );
  MX2X1 U789 ( .A(\iRF_stage/reg_bank/reg_bank[582] ), .B(n6), .S0(n616), .Y(
        \iRF_stage/reg_bank/n720 ) );
  MX2X1 U790 ( .A(\iRF_stage/reg_bank/reg_bank[581] ), .B(n7), .S0(n616), .Y(
        \iRF_stage/reg_bank/n719 ) );
  MX2X1 U791 ( .A(\iRF_stage/reg_bank/reg_bank[580] ), .B(n8), .S0(n616), .Y(
        \iRF_stage/reg_bank/n718 ) );
  MX2X1 U792 ( .A(\iRF_stage/reg_bank/reg_bank[579] ), .B(n9), .S0(n616), .Y(
        \iRF_stage/reg_bank/n717 ) );
  MX2X1 U793 ( .A(\iRF_stage/reg_bank/reg_bank[578] ), .B(n12), .S0(n616), .Y(
        \iRF_stage/reg_bank/n716 ) );
  MX2X1 U794 ( .A(\iRF_stage/reg_bank/reg_bank[577] ), .B(n23), .S0(n616), .Y(
        \iRF_stage/reg_bank/n715 ) );
  MX2X1 U795 ( .A(\iRF_stage/reg_bank/reg_bank[576] ), .B(n34), .S0(n616), .Y(
        \iRF_stage/reg_bank/n714 ) );
  AND2X1 U796 ( .A(n607), .B(n617), .Y(n616) );
  MX2X1 U797 ( .A(\iRF_stage/reg_bank/reg_bank[575] ), .B(n10), .S0(n618), .Y(
        \iRF_stage/reg_bank/n713 ) );
  MX2X1 U798 ( .A(\iRF_stage/reg_bank/reg_bank[574] ), .B(n11), .S0(n618), .Y(
        \iRF_stage/reg_bank/n712 ) );
  MX2X1 U799 ( .A(\iRF_stage/reg_bank/reg_bank[573] ), .B(n13), .S0(n618), .Y(
        \iRF_stage/reg_bank/n711 ) );
  MX2X1 U800 ( .A(\iRF_stage/reg_bank/reg_bank[572] ), .B(n14), .S0(n618), .Y(
        \iRF_stage/reg_bank/n710 ) );
  MX2X1 U801 ( .A(\iRF_stage/reg_bank/reg_bank[571] ), .B(n15), .S0(n618), .Y(
        \iRF_stage/reg_bank/n709 ) );
  MX2X1 U802 ( .A(\iRF_stage/reg_bank/reg_bank[570] ), .B(n16), .S0(n618), .Y(
        \iRF_stage/reg_bank/n708 ) );
  MX2X1 U803 ( .A(\iRF_stage/reg_bank/reg_bank[569] ), .B(n17), .S0(n618), .Y(
        \iRF_stage/reg_bank/n707 ) );
  MX2X1 U804 ( .A(\iRF_stage/reg_bank/reg_bank[568] ), .B(n18), .S0(n618), .Y(
        \iRF_stage/reg_bank/n706 ) );
  MX2X1 U805 ( .A(\iRF_stage/reg_bank/reg_bank[567] ), .B(n19), .S0(n618), .Y(
        \iRF_stage/reg_bank/n705 ) );
  MX2X1 U806 ( .A(\iRF_stage/reg_bank/reg_bank[566] ), .B(n20), .S0(n618), .Y(
        \iRF_stage/reg_bank/n704 ) );
  MX2X1 U807 ( .A(\iRF_stage/reg_bank/reg_bank[565] ), .B(n21), .S0(n618), .Y(
        \iRF_stage/reg_bank/n703 ) );
  MX2X1 U808 ( .A(\iRF_stage/reg_bank/reg_bank[564] ), .B(n22), .S0(n618), .Y(
        \iRF_stage/reg_bank/n702 ) );
  MX2X1 U809 ( .A(\iRF_stage/reg_bank/reg_bank[563] ), .B(n24), .S0(n618), .Y(
        \iRF_stage/reg_bank/n701 ) );
  MX2X1 U810 ( .A(\iRF_stage/reg_bank/reg_bank[562] ), .B(n25), .S0(n618), .Y(
        \iRF_stage/reg_bank/n700 ) );
  MX2X1 U811 ( .A(\iRF_stage/reg_bank/reg_bank[561] ), .B(n26), .S0(n618), .Y(
        \iRF_stage/reg_bank/n699 ) );
  MX2X1 U812 ( .A(\iRF_stage/reg_bank/reg_bank[560] ), .B(n27), .S0(n618), .Y(
        \iRF_stage/reg_bank/n698 ) );
  MX2X1 U813 ( .A(\iRF_stage/reg_bank/reg_bank[559] ), .B(n28), .S0(n618), .Y(
        \iRF_stage/reg_bank/n697 ) );
  MX2X1 U814 ( .A(\iRF_stage/reg_bank/reg_bank[558] ), .B(n29), .S0(n618), .Y(
        \iRF_stage/reg_bank/n696 ) );
  MX2X1 U815 ( .A(\iRF_stage/reg_bank/reg_bank[557] ), .B(n30), .S0(n618), .Y(
        \iRF_stage/reg_bank/n695 ) );
  MX2X1 U816 ( .A(\iRF_stage/reg_bank/reg_bank[556] ), .B(n31), .S0(n618), .Y(
        \iRF_stage/reg_bank/n694 ) );
  MX2X1 U817 ( .A(\iRF_stage/reg_bank/reg_bank[555] ), .B(n32), .S0(n618), .Y(
        \iRF_stage/reg_bank/n693 ) );
  MX2X1 U818 ( .A(\iRF_stage/reg_bank/reg_bank[554] ), .B(n33), .S0(n618), .Y(
        \iRF_stage/reg_bank/n692 ) );
  MX2X1 U819 ( .A(\iRF_stage/reg_bank/reg_bank[553] ), .B(n3), .S0(n618), .Y(
        \iRF_stage/reg_bank/n691 ) );
  MX2X1 U820 ( .A(\iRF_stage/reg_bank/reg_bank[552] ), .B(n4), .S0(n618), .Y(
        \iRF_stage/reg_bank/n690 ) );
  MX2X1 U821 ( .A(\iRF_stage/reg_bank/reg_bank[551] ), .B(n5), .S0(n618), .Y(
        \iRF_stage/reg_bank/n689 ) );
  MX2X1 U822 ( .A(\iRF_stage/reg_bank/reg_bank[550] ), .B(n6), .S0(n618), .Y(
        \iRF_stage/reg_bank/n688 ) );
  MX2X1 U823 ( .A(\iRF_stage/reg_bank/reg_bank[549] ), .B(n7), .S0(n618), .Y(
        \iRF_stage/reg_bank/n687 ) );
  MX2X1 U824 ( .A(\iRF_stage/reg_bank/reg_bank[548] ), .B(n8), .S0(n618), .Y(
        \iRF_stage/reg_bank/n686 ) );
  MX2X1 U825 ( .A(\iRF_stage/reg_bank/reg_bank[547] ), .B(n9), .S0(n618), .Y(
        \iRF_stage/reg_bank/n685 ) );
  MX2X1 U826 ( .A(\iRF_stage/reg_bank/reg_bank[546] ), .B(n12), .S0(n618), .Y(
        \iRF_stage/reg_bank/n684 ) );
  MX2X1 U827 ( .A(\iRF_stage/reg_bank/reg_bank[545] ), .B(n23), .S0(n618), .Y(
        \iRF_stage/reg_bank/n683 ) );
  MX2X1 U828 ( .A(\iRF_stage/reg_bank/reg_bank[544] ), .B(n34), .S0(n618), .Y(
        \iRF_stage/reg_bank/n682 ) );
  AND2X1 U829 ( .A(n607), .B(n601), .Y(n618) );
  MX2X1 U830 ( .A(\iRF_stage/reg_bank/reg_bank[543] ), .B(n10), .S0(n619), .Y(
        \iRF_stage/reg_bank/n681 ) );
  MX2X1 U831 ( .A(\iRF_stage/reg_bank/reg_bank[542] ), .B(n11), .S0(n619), .Y(
        \iRF_stage/reg_bank/n680 ) );
  MX2X1 U832 ( .A(\iRF_stage/reg_bank/reg_bank[541] ), .B(n13), .S0(n619), .Y(
        \iRF_stage/reg_bank/n679 ) );
  MX2X1 U833 ( .A(\iRF_stage/reg_bank/reg_bank[540] ), .B(n14), .S0(n619), .Y(
        \iRF_stage/reg_bank/n678 ) );
  MX2X1 U834 ( .A(\iRF_stage/reg_bank/reg_bank[539] ), .B(n15), .S0(n619), .Y(
        \iRF_stage/reg_bank/n677 ) );
  MX2X1 U835 ( .A(\iRF_stage/reg_bank/reg_bank[538] ), .B(n16), .S0(n619), .Y(
        \iRF_stage/reg_bank/n676 ) );
  MX2X1 U836 ( .A(\iRF_stage/reg_bank/reg_bank[537] ), .B(n17), .S0(n619), .Y(
        \iRF_stage/reg_bank/n675 ) );
  MX2X1 U837 ( .A(\iRF_stage/reg_bank/reg_bank[536] ), .B(n18), .S0(n619), .Y(
        \iRF_stage/reg_bank/n674 ) );
  MX2X1 U838 ( .A(\iRF_stage/reg_bank/reg_bank[535] ), .B(n19), .S0(n619), .Y(
        \iRF_stage/reg_bank/n673 ) );
  MX2X1 U839 ( .A(\iRF_stage/reg_bank/reg_bank[534] ), .B(n20), .S0(n619), .Y(
        \iRF_stage/reg_bank/n672 ) );
  MX2X1 U840 ( .A(\iRF_stage/reg_bank/reg_bank[533] ), .B(n21), .S0(n619), .Y(
        \iRF_stage/reg_bank/n671 ) );
  MX2X1 U841 ( .A(\iRF_stage/reg_bank/reg_bank[532] ), .B(n22), .S0(n619), .Y(
        \iRF_stage/reg_bank/n670 ) );
  MX2X1 U842 ( .A(\iRF_stage/reg_bank/reg_bank[531] ), .B(n24), .S0(n619), .Y(
        \iRF_stage/reg_bank/n669 ) );
  MX2X1 U843 ( .A(\iRF_stage/reg_bank/reg_bank[530] ), .B(n25), .S0(n619), .Y(
        \iRF_stage/reg_bank/n668 ) );
  MX2X1 U844 ( .A(\iRF_stage/reg_bank/reg_bank[529] ), .B(n26), .S0(n619), .Y(
        \iRF_stage/reg_bank/n667 ) );
  MX2X1 U845 ( .A(\iRF_stage/reg_bank/reg_bank[528] ), .B(n27), .S0(n619), .Y(
        \iRF_stage/reg_bank/n666 ) );
  MX2X1 U846 ( .A(\iRF_stage/reg_bank/reg_bank[527] ), .B(n28), .S0(n619), .Y(
        \iRF_stage/reg_bank/n665 ) );
  MX2X1 U847 ( .A(\iRF_stage/reg_bank/reg_bank[526] ), .B(n29), .S0(n619), .Y(
        \iRF_stage/reg_bank/n664 ) );
  MX2X1 U848 ( .A(\iRF_stage/reg_bank/reg_bank[525] ), .B(n30), .S0(n619), .Y(
        \iRF_stage/reg_bank/n663 ) );
  MX2X1 U849 ( .A(\iRF_stage/reg_bank/reg_bank[524] ), .B(n31), .S0(n619), .Y(
        \iRF_stage/reg_bank/n662 ) );
  MX2X1 U850 ( .A(\iRF_stage/reg_bank/reg_bank[523] ), .B(n32), .S0(n619), .Y(
        \iRF_stage/reg_bank/n661 ) );
  MX2X1 U851 ( .A(\iRF_stage/reg_bank/reg_bank[522] ), .B(n33), .S0(n619), .Y(
        \iRF_stage/reg_bank/n660 ) );
  MX2X1 U852 ( .A(\iRF_stage/reg_bank/reg_bank[521] ), .B(n3), .S0(n619), .Y(
        \iRF_stage/reg_bank/n659 ) );
  MX2X1 U853 ( .A(\iRF_stage/reg_bank/reg_bank[520] ), .B(n4), .S0(n619), .Y(
        \iRF_stage/reg_bank/n658 ) );
  MX2X1 U854 ( .A(\iRF_stage/reg_bank/reg_bank[519] ), .B(n5), .S0(n619), .Y(
        \iRF_stage/reg_bank/n657 ) );
  MX2X1 U855 ( .A(\iRF_stage/reg_bank/reg_bank[518] ), .B(n6), .S0(n619), .Y(
        \iRF_stage/reg_bank/n656 ) );
  MX2X1 U856 ( .A(\iRF_stage/reg_bank/reg_bank[517] ), .B(n7), .S0(n619), .Y(
        \iRF_stage/reg_bank/n655 ) );
  MX2X1 U857 ( .A(\iRF_stage/reg_bank/reg_bank[516] ), .B(n8), .S0(n619), .Y(
        \iRF_stage/reg_bank/n654 ) );
  MX2X1 U858 ( .A(\iRF_stage/reg_bank/reg_bank[515] ), .B(n9), .S0(n619), .Y(
        \iRF_stage/reg_bank/n653 ) );
  MX2X1 U859 ( .A(\iRF_stage/reg_bank/reg_bank[514] ), .B(n12), .S0(n619), .Y(
        \iRF_stage/reg_bank/n652 ) );
  MX2X1 U860 ( .A(\iRF_stage/reg_bank/reg_bank[513] ), .B(n23), .S0(n619), .Y(
        \iRF_stage/reg_bank/n651 ) );
  MX2X1 U861 ( .A(\iRF_stage/reg_bank/reg_bank[512] ), .B(n34), .S0(n619), .Y(
        \iRF_stage/reg_bank/n650 ) );
  AND2X1 U862 ( .A(n607), .B(n604), .Y(n619) );
  NOR3BX1 U863 ( .AN(\iRF_stage/reg_bank/r_wren ), .B(n620), .C(
        \iRF_stage/reg_bank/r_wraddress[4] ), .Y(n607) );
  MX2X1 U864 ( .A(\iRF_stage/reg_bank/reg_bank[511] ), .B(n10), .S0(n621), .Y(
        \iRF_stage/reg_bank/n649 ) );
  MX2X1 U865 ( .A(\iRF_stage/reg_bank/reg_bank[510] ), .B(n11), .S0(n621), .Y(
        \iRF_stage/reg_bank/n648 ) );
  MX2X1 U866 ( .A(\iRF_stage/reg_bank/reg_bank[509] ), .B(n13), .S0(n621), .Y(
        \iRF_stage/reg_bank/n647 ) );
  MX2X1 U867 ( .A(\iRF_stage/reg_bank/reg_bank[508] ), .B(n14), .S0(n621), .Y(
        \iRF_stage/reg_bank/n646 ) );
  MX2X1 U868 ( .A(\iRF_stage/reg_bank/reg_bank[507] ), .B(n15), .S0(n621), .Y(
        \iRF_stage/reg_bank/n645 ) );
  MX2X1 U869 ( .A(\iRF_stage/reg_bank/reg_bank[506] ), .B(n16), .S0(n621), .Y(
        \iRF_stage/reg_bank/n644 ) );
  MX2X1 U870 ( .A(\iRF_stage/reg_bank/reg_bank[505] ), .B(n17), .S0(n621), .Y(
        \iRF_stage/reg_bank/n643 ) );
  MX2X1 U871 ( .A(\iRF_stage/reg_bank/reg_bank[504] ), .B(n18), .S0(n621), .Y(
        \iRF_stage/reg_bank/n642 ) );
  MX2X1 U872 ( .A(\iRF_stage/reg_bank/reg_bank[503] ), .B(n19), .S0(n621), .Y(
        \iRF_stage/reg_bank/n641 ) );
  MX2X1 U873 ( .A(\iRF_stage/reg_bank/reg_bank[502] ), .B(n20), .S0(n621), .Y(
        \iRF_stage/reg_bank/n640 ) );
  MX2X1 U874 ( .A(\iRF_stage/reg_bank/reg_bank[501] ), .B(n21), .S0(n621), .Y(
        \iRF_stage/reg_bank/n639 ) );
  MX2X1 U875 ( .A(\iRF_stage/reg_bank/reg_bank[500] ), .B(n22), .S0(n621), .Y(
        \iRF_stage/reg_bank/n638 ) );
  MX2X1 U876 ( .A(\iRF_stage/reg_bank/reg_bank[499] ), .B(n24), .S0(n621), .Y(
        \iRF_stage/reg_bank/n637 ) );
  MX2X1 U877 ( .A(\iRF_stage/reg_bank/reg_bank[498] ), .B(n25), .S0(n621), .Y(
        \iRF_stage/reg_bank/n636 ) );
  MX2X1 U878 ( .A(\iRF_stage/reg_bank/reg_bank[497] ), .B(n26), .S0(n621), .Y(
        \iRF_stage/reg_bank/n635 ) );
  MX2X1 U879 ( .A(\iRF_stage/reg_bank/reg_bank[496] ), .B(n27), .S0(n621), .Y(
        \iRF_stage/reg_bank/n634 ) );
  MX2X1 U880 ( .A(\iRF_stage/reg_bank/reg_bank[495] ), .B(n28), .S0(n621), .Y(
        \iRF_stage/reg_bank/n633 ) );
  MX2X1 U881 ( .A(\iRF_stage/reg_bank/reg_bank[494] ), .B(n29), .S0(n621), .Y(
        \iRF_stage/reg_bank/n632 ) );
  MX2X1 U882 ( .A(\iRF_stage/reg_bank/reg_bank[493] ), .B(n30), .S0(n621), .Y(
        \iRF_stage/reg_bank/n631 ) );
  MX2X1 U883 ( .A(\iRF_stage/reg_bank/reg_bank[492] ), .B(n31), .S0(n621), .Y(
        \iRF_stage/reg_bank/n630 ) );
  MX2X1 U884 ( .A(\iRF_stage/reg_bank/reg_bank[491] ), .B(n32), .S0(n621), .Y(
        \iRF_stage/reg_bank/n629 ) );
  MX2X1 U885 ( .A(\iRF_stage/reg_bank/reg_bank[490] ), .B(n33), .S0(n621), .Y(
        \iRF_stage/reg_bank/n628 ) );
  MX2X1 U886 ( .A(\iRF_stage/reg_bank/reg_bank[489] ), .B(n3), .S0(n621), .Y(
        \iRF_stage/reg_bank/n627 ) );
  MX2X1 U887 ( .A(\iRF_stage/reg_bank/reg_bank[488] ), .B(n4), .S0(n621), .Y(
        \iRF_stage/reg_bank/n626 ) );
  MX2X1 U888 ( .A(\iRF_stage/reg_bank/reg_bank[487] ), .B(n5), .S0(n621), .Y(
        \iRF_stage/reg_bank/n625 ) );
  MX2X1 U889 ( .A(\iRF_stage/reg_bank/reg_bank[486] ), .B(n6), .S0(n621), .Y(
        \iRF_stage/reg_bank/n624 ) );
  MX2X1 U890 ( .A(\iRF_stage/reg_bank/reg_bank[485] ), .B(n7), .S0(n621), .Y(
        \iRF_stage/reg_bank/n623 ) );
  MX2X1 U891 ( .A(\iRF_stage/reg_bank/reg_bank[484] ), .B(n8), .S0(n621), .Y(
        \iRF_stage/reg_bank/n622 ) );
  MX2X1 U892 ( .A(\iRF_stage/reg_bank/reg_bank[483] ), .B(n9), .S0(n621), .Y(
        \iRF_stage/reg_bank/n621 ) );
  MX2X1 U893 ( .A(\iRF_stage/reg_bank/reg_bank[482] ), .B(n12), .S0(n621), .Y(
        \iRF_stage/reg_bank/n620 ) );
  MX2X1 U894 ( .A(\iRF_stage/reg_bank/reg_bank[481] ), .B(n23), .S0(n621), .Y(
        \iRF_stage/reg_bank/n619 ) );
  MX2X1 U895 ( .A(\iRF_stage/reg_bank/reg_bank[480] ), .B(n34), .S0(n621), .Y(
        \iRF_stage/reg_bank/n618 ) );
  AND2X1 U896 ( .A(n622), .B(n606), .Y(n621) );
  MX2X1 U897 ( .A(\iRF_stage/reg_bank/reg_bank[479] ), .B(n10), .S0(n623), .Y(
        \iRF_stage/reg_bank/n617 ) );
  MX2X1 U898 ( .A(\iRF_stage/reg_bank/reg_bank[478] ), .B(n11), .S0(n623), .Y(
        \iRF_stage/reg_bank/n616 ) );
  MX2X1 U899 ( .A(\iRF_stage/reg_bank/reg_bank[477] ), .B(n13), .S0(n623), .Y(
        \iRF_stage/reg_bank/n615 ) );
  MX2X1 U900 ( .A(\iRF_stage/reg_bank/reg_bank[476] ), .B(n14), .S0(n623), .Y(
        \iRF_stage/reg_bank/n614 ) );
  MX2X1 U901 ( .A(\iRF_stage/reg_bank/reg_bank[475] ), .B(n15), .S0(n623), .Y(
        \iRF_stage/reg_bank/n613 ) );
  MX2X1 U902 ( .A(\iRF_stage/reg_bank/reg_bank[474] ), .B(n16), .S0(n623), .Y(
        \iRF_stage/reg_bank/n612 ) );
  MX2X1 U903 ( .A(\iRF_stage/reg_bank/reg_bank[473] ), .B(n17), .S0(n623), .Y(
        \iRF_stage/reg_bank/n611 ) );
  MX2X1 U904 ( .A(\iRF_stage/reg_bank/reg_bank[472] ), .B(n18), .S0(n623), .Y(
        \iRF_stage/reg_bank/n610 ) );
  MX2X1 U905 ( .A(\iRF_stage/reg_bank/reg_bank[471] ), .B(n19), .S0(n623), .Y(
        \iRF_stage/reg_bank/n609 ) );
  MX2X1 U906 ( .A(\iRF_stage/reg_bank/reg_bank[470] ), .B(n20), .S0(n623), .Y(
        \iRF_stage/reg_bank/n608 ) );
  MX2X1 U907 ( .A(\iRF_stage/reg_bank/reg_bank[469] ), .B(n21), .S0(n623), .Y(
        \iRF_stage/reg_bank/n607 ) );
  MX2X1 U908 ( .A(\iRF_stage/reg_bank/reg_bank[468] ), .B(n22), .S0(n623), .Y(
        \iRF_stage/reg_bank/n606 ) );
  MX2X1 U909 ( .A(\iRF_stage/reg_bank/reg_bank[467] ), .B(n24), .S0(n623), .Y(
        \iRF_stage/reg_bank/n605 ) );
  MX2X1 U910 ( .A(\iRF_stage/reg_bank/reg_bank[466] ), .B(n25), .S0(n623), .Y(
        \iRF_stage/reg_bank/n604 ) );
  MX2X1 U911 ( .A(\iRF_stage/reg_bank/reg_bank[465] ), .B(n26), .S0(n623), .Y(
        \iRF_stage/reg_bank/n603 ) );
  MX2X1 U912 ( .A(\iRF_stage/reg_bank/reg_bank[464] ), .B(n27), .S0(n623), .Y(
        \iRF_stage/reg_bank/n602 ) );
  MX2X1 U913 ( .A(\iRF_stage/reg_bank/reg_bank[463] ), .B(n28), .S0(n623), .Y(
        \iRF_stage/reg_bank/n601 ) );
  MX2X1 U914 ( .A(\iRF_stage/reg_bank/reg_bank[462] ), .B(n29), .S0(n623), .Y(
        \iRF_stage/reg_bank/n600 ) );
  MX2X1 U915 ( .A(\iRF_stage/reg_bank/reg_bank[461] ), .B(n30), .S0(n623), .Y(
        \iRF_stage/reg_bank/n599 ) );
  MX2X1 U916 ( .A(\iRF_stage/reg_bank/reg_bank[460] ), .B(n31), .S0(n623), .Y(
        \iRF_stage/reg_bank/n598 ) );
  MX2X1 U917 ( .A(\iRF_stage/reg_bank/reg_bank[459] ), .B(n32), .S0(n623), .Y(
        \iRF_stage/reg_bank/n597 ) );
  MX2X1 U918 ( .A(\iRF_stage/reg_bank/reg_bank[458] ), .B(n33), .S0(n623), .Y(
        \iRF_stage/reg_bank/n596 ) );
  MX2X1 U919 ( .A(\iRF_stage/reg_bank/reg_bank[457] ), .B(n3), .S0(n623), .Y(
        \iRF_stage/reg_bank/n595 ) );
  MX2X1 U920 ( .A(\iRF_stage/reg_bank/reg_bank[456] ), .B(n4), .S0(n623), .Y(
        \iRF_stage/reg_bank/n594 ) );
  MX2X1 U921 ( .A(\iRF_stage/reg_bank/reg_bank[455] ), .B(n5), .S0(n623), .Y(
        \iRF_stage/reg_bank/n593 ) );
  MX2X1 U922 ( .A(\iRF_stage/reg_bank/reg_bank[454] ), .B(n6), .S0(n623), .Y(
        \iRF_stage/reg_bank/n592 ) );
  MX2X1 U923 ( .A(\iRF_stage/reg_bank/reg_bank[453] ), .B(n7), .S0(n623), .Y(
        \iRF_stage/reg_bank/n591 ) );
  MX2X1 U924 ( .A(\iRF_stage/reg_bank/reg_bank[452] ), .B(n8), .S0(n623), .Y(
        \iRF_stage/reg_bank/n590 ) );
  MX2X1 U925 ( .A(\iRF_stage/reg_bank/reg_bank[451] ), .B(n9), .S0(n623), .Y(
        \iRF_stage/reg_bank/n589 ) );
  MX2X1 U926 ( .A(\iRF_stage/reg_bank/reg_bank[450] ), .B(n12), .S0(n623), .Y(
        \iRF_stage/reg_bank/n588 ) );
  MX2X1 U927 ( .A(\iRF_stage/reg_bank/reg_bank[449] ), .B(n23), .S0(n623), .Y(
        \iRF_stage/reg_bank/n587 ) );
  MX2X1 U928 ( .A(\iRF_stage/reg_bank/reg_bank[448] ), .B(n34), .S0(n623), .Y(
        \iRF_stage/reg_bank/n586 ) );
  AND2X1 U929 ( .A(n622), .B(n609), .Y(n623) );
  MX2X1 U930 ( .A(\iRF_stage/reg_bank/reg_bank[447] ), .B(n10), .S0(n624), .Y(
        \iRF_stage/reg_bank/n585 ) );
  MX2X1 U931 ( .A(\iRF_stage/reg_bank/reg_bank[446] ), .B(n11), .S0(n624), .Y(
        \iRF_stage/reg_bank/n584 ) );
  MX2X1 U932 ( .A(\iRF_stage/reg_bank/reg_bank[445] ), .B(n13), .S0(n624), .Y(
        \iRF_stage/reg_bank/n583 ) );
  MX2X1 U933 ( .A(\iRF_stage/reg_bank/reg_bank[444] ), .B(n14), .S0(n624), .Y(
        \iRF_stage/reg_bank/n582 ) );
  MX2X1 U934 ( .A(\iRF_stage/reg_bank/reg_bank[443] ), .B(n15), .S0(n624), .Y(
        \iRF_stage/reg_bank/n581 ) );
  MX2X1 U935 ( .A(\iRF_stage/reg_bank/reg_bank[442] ), .B(n16), .S0(n624), .Y(
        \iRF_stage/reg_bank/n580 ) );
  MX2X1 U936 ( .A(\iRF_stage/reg_bank/reg_bank[441] ), .B(n17), .S0(n624), .Y(
        \iRF_stage/reg_bank/n579 ) );
  MX2X1 U937 ( .A(\iRF_stage/reg_bank/reg_bank[440] ), .B(n18), .S0(n624), .Y(
        \iRF_stage/reg_bank/n578 ) );
  MX2X1 U938 ( .A(\iRF_stage/reg_bank/reg_bank[439] ), .B(n19), .S0(n624), .Y(
        \iRF_stage/reg_bank/n577 ) );
  MX2X1 U939 ( .A(\iRF_stage/reg_bank/reg_bank[438] ), .B(n20), .S0(n624), .Y(
        \iRF_stage/reg_bank/n576 ) );
  MX2X1 U940 ( .A(\iRF_stage/reg_bank/reg_bank[437] ), .B(n21), .S0(n624), .Y(
        \iRF_stage/reg_bank/n575 ) );
  MX2X1 U941 ( .A(\iRF_stage/reg_bank/reg_bank[436] ), .B(n22), .S0(n624), .Y(
        \iRF_stage/reg_bank/n574 ) );
  MX2X1 U942 ( .A(\iRF_stage/reg_bank/reg_bank[435] ), .B(n24), .S0(n624), .Y(
        \iRF_stage/reg_bank/n573 ) );
  MX2X1 U943 ( .A(\iRF_stage/reg_bank/reg_bank[434] ), .B(n25), .S0(n624), .Y(
        \iRF_stage/reg_bank/n572 ) );
  MX2X1 U944 ( .A(\iRF_stage/reg_bank/reg_bank[433] ), .B(n26), .S0(n624), .Y(
        \iRF_stage/reg_bank/n571 ) );
  MX2X1 U945 ( .A(\iRF_stage/reg_bank/reg_bank[432] ), .B(n27), .S0(n624), .Y(
        \iRF_stage/reg_bank/n570 ) );
  MX2X1 U946 ( .A(\iRF_stage/reg_bank/reg_bank[431] ), .B(n28), .S0(n624), .Y(
        \iRF_stage/reg_bank/n569 ) );
  MX2X1 U947 ( .A(\iRF_stage/reg_bank/reg_bank[430] ), .B(n29), .S0(n624), .Y(
        \iRF_stage/reg_bank/n568 ) );
  MX2X1 U948 ( .A(\iRF_stage/reg_bank/reg_bank[429] ), .B(n30), .S0(n624), .Y(
        \iRF_stage/reg_bank/n567 ) );
  MX2X1 U949 ( .A(\iRF_stage/reg_bank/reg_bank[428] ), .B(n31), .S0(n624), .Y(
        \iRF_stage/reg_bank/n566 ) );
  MX2X1 U950 ( .A(\iRF_stage/reg_bank/reg_bank[427] ), .B(n32), .S0(n624), .Y(
        \iRF_stage/reg_bank/n565 ) );
  MX2X1 U951 ( .A(\iRF_stage/reg_bank/reg_bank[426] ), .B(n33), .S0(n624), .Y(
        \iRF_stage/reg_bank/n564 ) );
  MX2X1 U952 ( .A(\iRF_stage/reg_bank/reg_bank[425] ), .B(n3), .S0(n624), .Y(
        \iRF_stage/reg_bank/n563 ) );
  MX2X1 U953 ( .A(\iRF_stage/reg_bank/reg_bank[424] ), .B(n4), .S0(n624), .Y(
        \iRF_stage/reg_bank/n562 ) );
  MX2X1 U954 ( .A(\iRF_stage/reg_bank/reg_bank[423] ), .B(n5), .S0(n624), .Y(
        \iRF_stage/reg_bank/n561 ) );
  MX2X1 U955 ( .A(\iRF_stage/reg_bank/reg_bank[422] ), .B(n6), .S0(n624), .Y(
        \iRF_stage/reg_bank/n560 ) );
  MX2X1 U956 ( .A(\iRF_stage/reg_bank/reg_bank[421] ), .B(n7), .S0(n624), .Y(
        \iRF_stage/reg_bank/n559 ) );
  MX2X1 U957 ( .A(\iRF_stage/reg_bank/reg_bank[420] ), .B(n8), .S0(n624), .Y(
        \iRF_stage/reg_bank/n558 ) );
  MX2X1 U958 ( .A(\iRF_stage/reg_bank/reg_bank[419] ), .B(n9), .S0(n624), .Y(
        \iRF_stage/reg_bank/n557 ) );
  MX2X1 U959 ( .A(\iRF_stage/reg_bank/reg_bank[418] ), .B(n12), .S0(n624), .Y(
        \iRF_stage/reg_bank/n556 ) );
  MX2X1 U960 ( .A(\iRF_stage/reg_bank/reg_bank[417] ), .B(n23), .S0(n624), .Y(
        \iRF_stage/reg_bank/n555 ) );
  MX2X1 U961 ( .A(\iRF_stage/reg_bank/reg_bank[416] ), .B(n34), .S0(n624), .Y(
        \iRF_stage/reg_bank/n554 ) );
  AND2X1 U962 ( .A(n622), .B(n611), .Y(n624) );
  MX2X1 U963 ( .A(\iRF_stage/reg_bank/reg_bank[415] ), .B(n10), .S0(n625), .Y(
        \iRF_stage/reg_bank/n553 ) );
  MX2X1 U964 ( .A(\iRF_stage/reg_bank/reg_bank[414] ), .B(n11), .S0(n625), .Y(
        \iRF_stage/reg_bank/n552 ) );
  MX2X1 U965 ( .A(\iRF_stage/reg_bank/reg_bank[413] ), .B(n13), .S0(n625), .Y(
        \iRF_stage/reg_bank/n551 ) );
  MX2X1 U966 ( .A(\iRF_stage/reg_bank/reg_bank[412] ), .B(n14), .S0(n625), .Y(
        \iRF_stage/reg_bank/n550 ) );
  MX2X1 U967 ( .A(\iRF_stage/reg_bank/reg_bank[411] ), .B(n15), .S0(n625), .Y(
        \iRF_stage/reg_bank/n549 ) );
  MX2X1 U968 ( .A(\iRF_stage/reg_bank/reg_bank[410] ), .B(n16), .S0(n625), .Y(
        \iRF_stage/reg_bank/n548 ) );
  MX2X1 U969 ( .A(\iRF_stage/reg_bank/reg_bank[409] ), .B(n17), .S0(n625), .Y(
        \iRF_stage/reg_bank/n547 ) );
  MX2X1 U970 ( .A(\iRF_stage/reg_bank/reg_bank[408] ), .B(n18), .S0(n625), .Y(
        \iRF_stage/reg_bank/n546 ) );
  MX2X1 U971 ( .A(\iRF_stage/reg_bank/reg_bank[407] ), .B(n19), .S0(n625), .Y(
        \iRF_stage/reg_bank/n545 ) );
  MX2X1 U972 ( .A(\iRF_stage/reg_bank/reg_bank[406] ), .B(n20), .S0(n625), .Y(
        \iRF_stage/reg_bank/n544 ) );
  MX2X1 U973 ( .A(\iRF_stage/reg_bank/reg_bank[405] ), .B(n21), .S0(n625), .Y(
        \iRF_stage/reg_bank/n543 ) );
  MX2X1 U974 ( .A(\iRF_stage/reg_bank/reg_bank[404] ), .B(n22), .S0(n625), .Y(
        \iRF_stage/reg_bank/n542 ) );
  MX2X1 U975 ( .A(\iRF_stage/reg_bank/reg_bank[403] ), .B(n24), .S0(n625), .Y(
        \iRF_stage/reg_bank/n541 ) );
  MX2X1 U976 ( .A(\iRF_stage/reg_bank/reg_bank[402] ), .B(n25), .S0(n625), .Y(
        \iRF_stage/reg_bank/n540 ) );
  MX2X1 U977 ( .A(\iRF_stage/reg_bank/reg_bank[401] ), .B(n26), .S0(n625), .Y(
        \iRF_stage/reg_bank/n539 ) );
  MX2X1 U978 ( .A(\iRF_stage/reg_bank/reg_bank[400] ), .B(n27), .S0(n625), .Y(
        \iRF_stage/reg_bank/n538 ) );
  MX2X1 U979 ( .A(\iRF_stage/reg_bank/reg_bank[399] ), .B(n28), .S0(n625), .Y(
        \iRF_stage/reg_bank/n537 ) );
  MX2X1 U980 ( .A(\iRF_stage/reg_bank/reg_bank[398] ), .B(n29), .S0(n625), .Y(
        \iRF_stage/reg_bank/n536 ) );
  MX2X1 U981 ( .A(\iRF_stage/reg_bank/reg_bank[397] ), .B(n30), .S0(n625), .Y(
        \iRF_stage/reg_bank/n535 ) );
  MX2X1 U982 ( .A(\iRF_stage/reg_bank/reg_bank[396] ), .B(n31), .S0(n625), .Y(
        \iRF_stage/reg_bank/n534 ) );
  MX2X1 U983 ( .A(\iRF_stage/reg_bank/reg_bank[395] ), .B(n32), .S0(n625), .Y(
        \iRF_stage/reg_bank/n533 ) );
  MX2X1 U984 ( .A(\iRF_stage/reg_bank/reg_bank[394] ), .B(n33), .S0(n625), .Y(
        \iRF_stage/reg_bank/n532 ) );
  MX2X1 U985 ( .A(\iRF_stage/reg_bank/reg_bank[393] ), .B(n3), .S0(n625), .Y(
        \iRF_stage/reg_bank/n531 ) );
  MX2X1 U986 ( .A(\iRF_stage/reg_bank/reg_bank[392] ), .B(n4), .S0(n625), .Y(
        \iRF_stage/reg_bank/n530 ) );
  MX2X1 U987 ( .A(\iRF_stage/reg_bank/reg_bank[391] ), .B(n5), .S0(n625), .Y(
        \iRF_stage/reg_bank/n529 ) );
  MX2X1 U988 ( .A(\iRF_stage/reg_bank/reg_bank[390] ), .B(n6), .S0(n625), .Y(
        \iRF_stage/reg_bank/n528 ) );
  MX2X1 U989 ( .A(\iRF_stage/reg_bank/reg_bank[389] ), .B(n7), .S0(n625), .Y(
        \iRF_stage/reg_bank/n527 ) );
  MX2X1 U990 ( .A(\iRF_stage/reg_bank/reg_bank[388] ), .B(n8), .S0(n625), .Y(
        \iRF_stage/reg_bank/n526 ) );
  MX2X1 U991 ( .A(\iRF_stage/reg_bank/reg_bank[387] ), .B(n9), .S0(n625), .Y(
        \iRF_stage/reg_bank/n525 ) );
  MX2X1 U992 ( .A(\iRF_stage/reg_bank/reg_bank[386] ), .B(n12), .S0(n625), .Y(
        \iRF_stage/reg_bank/n524 ) );
  MX2X1 U993 ( .A(\iRF_stage/reg_bank/reg_bank[385] ), .B(n23), .S0(n625), .Y(
        \iRF_stage/reg_bank/n523 ) );
  MX2X1 U994 ( .A(\iRF_stage/reg_bank/reg_bank[384] ), .B(n34), .S0(n625), .Y(
        \iRF_stage/reg_bank/n522 ) );
  AND2X1 U995 ( .A(n622), .B(n613), .Y(n625) );
  MX2X1 U996 ( .A(\iRF_stage/reg_bank/reg_bank[383] ), .B(n10), .S0(n626), .Y(
        \iRF_stage/reg_bank/n521 ) );
  MX2X1 U997 ( .A(\iRF_stage/reg_bank/reg_bank[382] ), .B(n11), .S0(n626), .Y(
        \iRF_stage/reg_bank/n520 ) );
  MX2X1 U998 ( .A(\iRF_stage/reg_bank/reg_bank[381] ), .B(n13), .S0(n626), .Y(
        \iRF_stage/reg_bank/n519 ) );
  MX2X1 U999 ( .A(\iRF_stage/reg_bank/reg_bank[380] ), .B(n14), .S0(n626), .Y(
        \iRF_stage/reg_bank/n518 ) );
  MX2X1 U1000 ( .A(\iRF_stage/reg_bank/reg_bank[379] ), .B(n15), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n517 ) );
  MX2X1 U1001 ( .A(\iRF_stage/reg_bank/reg_bank[378] ), .B(n16), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n516 ) );
  MX2X1 U1002 ( .A(\iRF_stage/reg_bank/reg_bank[377] ), .B(n17), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n515 ) );
  MX2X1 U1003 ( .A(\iRF_stage/reg_bank/reg_bank[376] ), .B(n18), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n514 ) );
  MX2X1 U1004 ( .A(\iRF_stage/reg_bank/reg_bank[375] ), .B(n19), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n513 ) );
  MX2X1 U1005 ( .A(\iRF_stage/reg_bank/reg_bank[374] ), .B(n20), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n512 ) );
  MX2X1 U1006 ( .A(\iRF_stage/reg_bank/reg_bank[373] ), .B(n21), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n511 ) );
  MX2X1 U1007 ( .A(\iRF_stage/reg_bank/reg_bank[372] ), .B(n22), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n510 ) );
  MX2X1 U1008 ( .A(\iRF_stage/reg_bank/reg_bank[371] ), .B(n24), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n509 ) );
  MX2X1 U1009 ( .A(\iRF_stage/reg_bank/reg_bank[370] ), .B(n25), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n508 ) );
  MX2X1 U1010 ( .A(\iRF_stage/reg_bank/reg_bank[369] ), .B(n26), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n507 ) );
  MX2X1 U1011 ( .A(\iRF_stage/reg_bank/reg_bank[368] ), .B(n27), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n506 ) );
  MX2X1 U1012 ( .A(\iRF_stage/reg_bank/reg_bank[367] ), .B(n28), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n505 ) );
  MX2X1 U1013 ( .A(\iRF_stage/reg_bank/reg_bank[366] ), .B(n29), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n504 ) );
  MX2X1 U1014 ( .A(\iRF_stage/reg_bank/reg_bank[365] ), .B(n30), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n503 ) );
  MX2X1 U1015 ( .A(\iRF_stage/reg_bank/reg_bank[364] ), .B(n31), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n502 ) );
  MX2X1 U1016 ( .A(\iRF_stage/reg_bank/reg_bank[363] ), .B(n32), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n501 ) );
  MX2X1 U1017 ( .A(\iRF_stage/reg_bank/reg_bank[362] ), .B(n33), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n500 ) );
  MX2X1 U1018 ( .A(\iRF_stage/reg_bank/reg_bank[361] ), .B(n3), .S0(n626), .Y(
        \iRF_stage/reg_bank/n499 ) );
  MX2X1 U1019 ( .A(\iRF_stage/reg_bank/reg_bank[360] ), .B(n4), .S0(n626), .Y(
        \iRF_stage/reg_bank/n498 ) );
  MX2X1 U1020 ( .A(\iRF_stage/reg_bank/reg_bank[359] ), .B(n5), .S0(n626), .Y(
        \iRF_stage/reg_bank/n497 ) );
  MX2X1 U1021 ( .A(\iRF_stage/reg_bank/reg_bank[358] ), .B(n6), .S0(n626), .Y(
        \iRF_stage/reg_bank/n496 ) );
  MX2X1 U1022 ( .A(\iRF_stage/reg_bank/reg_bank[357] ), .B(n7), .S0(n626), .Y(
        \iRF_stage/reg_bank/n495 ) );
  MX2X1 U1023 ( .A(\iRF_stage/reg_bank/reg_bank[356] ), .B(n8), .S0(n626), .Y(
        \iRF_stage/reg_bank/n494 ) );
  MX2X1 U1024 ( .A(\iRF_stage/reg_bank/reg_bank[355] ), .B(n9), .S0(n626), .Y(
        \iRF_stage/reg_bank/n493 ) );
  MX2X1 U1025 ( .A(\iRF_stage/reg_bank/reg_bank[354] ), .B(n12), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n492 ) );
  MX2X1 U1026 ( .A(\iRF_stage/reg_bank/reg_bank[353] ), .B(n23), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n491 ) );
  MX2X1 U1027 ( .A(\iRF_stage/reg_bank/reg_bank[352] ), .B(n34), .S0(n626), 
        .Y(\iRF_stage/reg_bank/n490 ) );
  AND2X1 U1028 ( .A(n622), .B(n615), .Y(n626) );
  MX2X1 U1029 ( .A(\iRF_stage/reg_bank/reg_bank[351] ), .B(n10), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n489 ) );
  MX2X1 U1030 ( .A(\iRF_stage/reg_bank/reg_bank[350] ), .B(n11), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n488 ) );
  MX2X1 U1031 ( .A(\iRF_stage/reg_bank/reg_bank[349] ), .B(n13), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n487 ) );
  MX2X1 U1032 ( .A(\iRF_stage/reg_bank/reg_bank[348] ), .B(n14), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n486 ) );
  MX2X1 U1033 ( .A(\iRF_stage/reg_bank/reg_bank[347] ), .B(n15), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n485 ) );
  MX2X1 U1034 ( .A(\iRF_stage/reg_bank/reg_bank[346] ), .B(n16), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n484 ) );
  MX2X1 U1035 ( .A(\iRF_stage/reg_bank/reg_bank[345] ), .B(n17), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n483 ) );
  MX2X1 U1036 ( .A(\iRF_stage/reg_bank/reg_bank[344] ), .B(n18), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n482 ) );
  MX2X1 U1037 ( .A(\iRF_stage/reg_bank/reg_bank[343] ), .B(n19), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n481 ) );
  MX2X1 U1038 ( .A(\iRF_stage/reg_bank/reg_bank[342] ), .B(n20), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n480 ) );
  MX2X1 U1039 ( .A(\iRF_stage/reg_bank/reg_bank[341] ), .B(n21), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n479 ) );
  MX2X1 U1040 ( .A(\iRF_stage/reg_bank/reg_bank[340] ), .B(n22), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n478 ) );
  MX2X1 U1041 ( .A(\iRF_stage/reg_bank/reg_bank[339] ), .B(n24), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n477 ) );
  MX2X1 U1042 ( .A(\iRF_stage/reg_bank/reg_bank[338] ), .B(n25), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n476 ) );
  MX2X1 U1043 ( .A(\iRF_stage/reg_bank/reg_bank[337] ), .B(n26), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n475 ) );
  MX2X1 U1044 ( .A(\iRF_stage/reg_bank/reg_bank[336] ), .B(n27), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n474 ) );
  MX2X1 U1045 ( .A(\iRF_stage/reg_bank/reg_bank[335] ), .B(n28), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n473 ) );
  MX2X1 U1046 ( .A(\iRF_stage/reg_bank/reg_bank[334] ), .B(n29), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n472 ) );
  MX2X1 U1047 ( .A(\iRF_stage/reg_bank/reg_bank[333] ), .B(n30), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n471 ) );
  MX2X1 U1048 ( .A(\iRF_stage/reg_bank/reg_bank[332] ), .B(n31), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n470 ) );
  MX2X1 U1049 ( .A(\iRF_stage/reg_bank/reg_bank[331] ), .B(n32), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n469 ) );
  MX2X1 U1050 ( .A(\iRF_stage/reg_bank/reg_bank[330] ), .B(n33), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n468 ) );
  MX2X1 U1051 ( .A(\iRF_stage/reg_bank/reg_bank[329] ), .B(n3), .S0(n627), .Y(
        \iRF_stage/reg_bank/n467 ) );
  MX2X1 U1052 ( .A(\iRF_stage/reg_bank/reg_bank[328] ), .B(n4), .S0(n627), .Y(
        \iRF_stage/reg_bank/n466 ) );
  MX2X1 U1053 ( .A(\iRF_stage/reg_bank/reg_bank[327] ), .B(n5), .S0(n627), .Y(
        \iRF_stage/reg_bank/n465 ) );
  MX2X1 U1054 ( .A(\iRF_stage/reg_bank/reg_bank[326] ), .B(n6), .S0(n627), .Y(
        \iRF_stage/reg_bank/n464 ) );
  MX2X1 U1055 ( .A(\iRF_stage/reg_bank/reg_bank[325] ), .B(n7), .S0(n627), .Y(
        \iRF_stage/reg_bank/n463 ) );
  MX2X1 U1056 ( .A(\iRF_stage/reg_bank/reg_bank[324] ), .B(n8), .S0(n627), .Y(
        \iRF_stage/reg_bank/n462 ) );
  MX2X1 U1057 ( .A(\iRF_stage/reg_bank/reg_bank[323] ), .B(n9), .S0(n627), .Y(
        \iRF_stage/reg_bank/n461 ) );
  MX2X1 U1058 ( .A(\iRF_stage/reg_bank/reg_bank[322] ), .B(n12), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n460 ) );
  MX2X1 U1059 ( .A(\iRF_stage/reg_bank/reg_bank[321] ), .B(n23), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n459 ) );
  MX2X1 U1060 ( .A(\iRF_stage/reg_bank/reg_bank[320] ), .B(n34), .S0(n627), 
        .Y(\iRF_stage/reg_bank/n458 ) );
  AND2X1 U1061 ( .A(n622), .B(n617), .Y(n627) );
  MX2X1 U1062 ( .A(\iRF_stage/reg_bank/reg_bank[319] ), .B(n10), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n457 ) );
  MX2X1 U1063 ( .A(\iRF_stage/reg_bank/reg_bank[318] ), .B(n11), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n456 ) );
  MX2X1 U1064 ( .A(\iRF_stage/reg_bank/reg_bank[317] ), .B(n13), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n455 ) );
  MX2X1 U1065 ( .A(\iRF_stage/reg_bank/reg_bank[316] ), .B(n14), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n454 ) );
  MX2X1 U1066 ( .A(\iRF_stage/reg_bank/reg_bank[315] ), .B(n15), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n453 ) );
  MX2X1 U1067 ( .A(\iRF_stage/reg_bank/reg_bank[314] ), .B(n16), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n452 ) );
  MX2X1 U1068 ( .A(\iRF_stage/reg_bank/reg_bank[313] ), .B(n17), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n451 ) );
  MX2X1 U1069 ( .A(\iRF_stage/reg_bank/reg_bank[312] ), .B(n18), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n450 ) );
  MX2X1 U1070 ( .A(\iRF_stage/reg_bank/reg_bank[311] ), .B(n19), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n449 ) );
  MX2X1 U1071 ( .A(\iRF_stage/reg_bank/reg_bank[310] ), .B(n20), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n448 ) );
  MX2X1 U1072 ( .A(\iRF_stage/reg_bank/reg_bank[309] ), .B(n21), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n447 ) );
  MX2X1 U1073 ( .A(\iRF_stage/reg_bank/reg_bank[308] ), .B(n22), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n446 ) );
  MX2X1 U1074 ( .A(\iRF_stage/reg_bank/reg_bank[307] ), .B(n24), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n445 ) );
  MX2X1 U1075 ( .A(\iRF_stage/reg_bank/reg_bank[306] ), .B(n25), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n444 ) );
  MX2X1 U1076 ( .A(\iRF_stage/reg_bank/reg_bank[305] ), .B(n26), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n443 ) );
  MX2X1 U1077 ( .A(\iRF_stage/reg_bank/reg_bank[304] ), .B(n27), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n442 ) );
  MX2X1 U1078 ( .A(\iRF_stage/reg_bank/reg_bank[303] ), .B(n28), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n441 ) );
  MX2X1 U1079 ( .A(\iRF_stage/reg_bank/reg_bank[302] ), .B(n29), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n440 ) );
  MX2X1 U1080 ( .A(\iRF_stage/reg_bank/reg_bank[301] ), .B(n30), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n439 ) );
  MX2X1 U1081 ( .A(\iRF_stage/reg_bank/reg_bank[300] ), .B(n31), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n438 ) );
  MX2X1 U1082 ( .A(\iRF_stage/reg_bank/reg_bank[299] ), .B(n32), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n437 ) );
  MX2X1 U1083 ( .A(\iRF_stage/reg_bank/reg_bank[298] ), .B(n33), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n436 ) );
  MX2X1 U1084 ( .A(\iRF_stage/reg_bank/reg_bank[297] ), .B(n3), .S0(n628), .Y(
        \iRF_stage/reg_bank/n435 ) );
  MX2X1 U1085 ( .A(\iRF_stage/reg_bank/reg_bank[296] ), .B(n4), .S0(n628), .Y(
        \iRF_stage/reg_bank/n434 ) );
  MX2X1 U1086 ( .A(\iRF_stage/reg_bank/reg_bank[295] ), .B(n5), .S0(n628), .Y(
        \iRF_stage/reg_bank/n433 ) );
  MX2X1 U1087 ( .A(\iRF_stage/reg_bank/reg_bank[294] ), .B(n6), .S0(n628), .Y(
        \iRF_stage/reg_bank/n432 ) );
  MX2X1 U1088 ( .A(\iRF_stage/reg_bank/reg_bank[293] ), .B(n7), .S0(n628), .Y(
        \iRF_stage/reg_bank/n431 ) );
  MX2X1 U1089 ( .A(\iRF_stage/reg_bank/reg_bank[292] ), .B(n8), .S0(n628), .Y(
        \iRF_stage/reg_bank/n430 ) );
  MX2X1 U1090 ( .A(\iRF_stage/reg_bank/reg_bank[291] ), .B(n9), .S0(n628), .Y(
        \iRF_stage/reg_bank/n429 ) );
  MX2X1 U1091 ( .A(\iRF_stage/reg_bank/reg_bank[290] ), .B(n12), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n428 ) );
  MX2X1 U1092 ( .A(\iRF_stage/reg_bank/reg_bank[289] ), .B(n23), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n427 ) );
  MX2X1 U1093 ( .A(\iRF_stage/reg_bank/reg_bank[288] ), .B(n34), .S0(n628), 
        .Y(\iRF_stage/reg_bank/n426 ) );
  AND2X1 U1094 ( .A(n622), .B(n601), .Y(n628) );
  MX2X1 U1095 ( .A(\iRF_stage/reg_bank/reg_bank[287] ), .B(n10), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n425 ) );
  MX2X1 U1096 ( .A(\iRF_stage/reg_bank/reg_bank[286] ), .B(n11), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n424 ) );
  MX2X1 U1097 ( .A(\iRF_stage/reg_bank/reg_bank[285] ), .B(n13), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n423 ) );
  MX2X1 U1098 ( .A(\iRF_stage/reg_bank/reg_bank[284] ), .B(n14), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n422 ) );
  MX2X1 U1099 ( .A(\iRF_stage/reg_bank/reg_bank[283] ), .B(n15), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n421 ) );
  MX2X1 U1100 ( .A(\iRF_stage/reg_bank/reg_bank[282] ), .B(n16), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n420 ) );
  MX2X1 U1101 ( .A(\iRF_stage/reg_bank/reg_bank[281] ), .B(n17), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n419 ) );
  MX2X1 U1102 ( .A(\iRF_stage/reg_bank/reg_bank[280] ), .B(n18), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n418 ) );
  MX2X1 U1103 ( .A(\iRF_stage/reg_bank/reg_bank[279] ), .B(n19), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n417 ) );
  MX2X1 U1104 ( .A(\iRF_stage/reg_bank/reg_bank[278] ), .B(n20), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n416 ) );
  MX2X1 U1105 ( .A(\iRF_stage/reg_bank/reg_bank[277] ), .B(n21), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n415 ) );
  MX2X1 U1106 ( .A(\iRF_stage/reg_bank/reg_bank[276] ), .B(n22), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n414 ) );
  MX2X1 U1107 ( .A(\iRF_stage/reg_bank/reg_bank[275] ), .B(n24), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n413 ) );
  MX2X1 U1108 ( .A(\iRF_stage/reg_bank/reg_bank[274] ), .B(n25), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n412 ) );
  MX2X1 U1109 ( .A(\iRF_stage/reg_bank/reg_bank[273] ), .B(n26), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n411 ) );
  MX2X1 U1110 ( .A(\iRF_stage/reg_bank/reg_bank[272] ), .B(n27), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n410 ) );
  MX2X1 U1111 ( .A(\iRF_stage/reg_bank/reg_bank[271] ), .B(n28), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n409 ) );
  MX2X1 U1112 ( .A(\iRF_stage/reg_bank/reg_bank[270] ), .B(n29), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n408 ) );
  MX2X1 U1113 ( .A(\iRF_stage/reg_bank/reg_bank[269] ), .B(n30), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n407 ) );
  MX2X1 U1114 ( .A(\iRF_stage/reg_bank/reg_bank[268] ), .B(n31), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n406 ) );
  MX2X1 U1115 ( .A(\iRF_stage/reg_bank/reg_bank[267] ), .B(n32), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n405 ) );
  MX2X1 U1116 ( .A(\iRF_stage/reg_bank/reg_bank[266] ), .B(n33), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n404 ) );
  MX2X1 U1117 ( .A(\iRF_stage/reg_bank/reg_bank[265] ), .B(n3), .S0(n629), .Y(
        \iRF_stage/reg_bank/n403 ) );
  MX2X1 U1118 ( .A(\iRF_stage/reg_bank/reg_bank[264] ), .B(n4), .S0(n629), .Y(
        \iRF_stage/reg_bank/n402 ) );
  MX2X1 U1119 ( .A(\iRF_stage/reg_bank/reg_bank[263] ), .B(n5), .S0(n629), .Y(
        \iRF_stage/reg_bank/n401 ) );
  MX2X1 U1120 ( .A(\iRF_stage/reg_bank/reg_bank[262] ), .B(n6), .S0(n629), .Y(
        \iRF_stage/reg_bank/n400 ) );
  MX2X1 U1121 ( .A(\iRF_stage/reg_bank/reg_bank[261] ), .B(n7), .S0(n629), .Y(
        \iRF_stage/reg_bank/n399 ) );
  MX2X1 U1122 ( .A(\iRF_stage/reg_bank/reg_bank[260] ), .B(n8), .S0(n629), .Y(
        \iRF_stage/reg_bank/n398 ) );
  MX2X1 U1123 ( .A(\iRF_stage/reg_bank/reg_bank[259] ), .B(n9), .S0(n629), .Y(
        \iRF_stage/reg_bank/n397 ) );
  MX2X1 U1124 ( .A(\iRF_stage/reg_bank/reg_bank[258] ), .B(n12), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n396 ) );
  MX2X1 U1125 ( .A(\iRF_stage/reg_bank/reg_bank[257] ), .B(n23), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n395 ) );
  MX2X1 U1126 ( .A(\iRF_stage/reg_bank/reg_bank[256] ), .B(n34), .S0(n629), 
        .Y(\iRF_stage/reg_bank/n394 ) );
  AND2X1 U1127 ( .A(n622), .B(n604), .Y(n629) );
  NOR3BX1 U1128 ( .AN(\iRF_stage/reg_bank/r_wren ), .B(n630), .C(
        \iRF_stage/reg_bank/r_wraddress[3] ), .Y(n622) );
  MX2X1 U1129 ( .A(\iRF_stage/reg_bank/reg_bank[255] ), .B(n10), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n393 ) );
  MX2X1 U1130 ( .A(\iRF_stage/reg_bank/reg_bank[254] ), .B(n11), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n392 ) );
  MX2X1 U1131 ( .A(\iRF_stage/reg_bank/reg_bank[253] ), .B(n13), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n391 ) );
  MX2X1 U1132 ( .A(\iRF_stage/reg_bank/reg_bank[252] ), .B(n14), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n390 ) );
  MX2X1 U1133 ( .A(\iRF_stage/reg_bank/reg_bank[251] ), .B(n15), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n389 ) );
  MX2X1 U1134 ( .A(\iRF_stage/reg_bank/reg_bank[250] ), .B(n16), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n388 ) );
  MX2X1 U1135 ( .A(\iRF_stage/reg_bank/reg_bank[249] ), .B(n17), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n387 ) );
  MX2X1 U1136 ( .A(\iRF_stage/reg_bank/reg_bank[248] ), .B(n18), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n386 ) );
  MX2X1 U1137 ( .A(\iRF_stage/reg_bank/reg_bank[247] ), .B(n19), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n385 ) );
  MX2X1 U1138 ( .A(\iRF_stage/reg_bank/reg_bank[246] ), .B(n20), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n384 ) );
  MX2X1 U1139 ( .A(\iRF_stage/reg_bank/reg_bank[245] ), .B(n21), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n383 ) );
  MX2X1 U1140 ( .A(\iRF_stage/reg_bank/reg_bank[244] ), .B(n22), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n382 ) );
  MX2X1 U1141 ( .A(\iRF_stage/reg_bank/reg_bank[243] ), .B(n24), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n381 ) );
  MX2X1 U1142 ( .A(\iRF_stage/reg_bank/reg_bank[242] ), .B(n25), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n380 ) );
  MX2X1 U1143 ( .A(\iRF_stage/reg_bank/reg_bank[241] ), .B(n26), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n379 ) );
  MX2X1 U1144 ( .A(\iRF_stage/reg_bank/reg_bank[240] ), .B(n27), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n378 ) );
  MX2X1 U1145 ( .A(\iRF_stage/reg_bank/reg_bank[239] ), .B(n28), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n377 ) );
  MX2X1 U1146 ( .A(\iRF_stage/reg_bank/reg_bank[238] ), .B(n29), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n376 ) );
  MX2X1 U1147 ( .A(\iRF_stage/reg_bank/reg_bank[237] ), .B(n30), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n375 ) );
  MX2X1 U1148 ( .A(\iRF_stage/reg_bank/reg_bank[236] ), .B(n31), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n374 ) );
  MX2X1 U1149 ( .A(\iRF_stage/reg_bank/reg_bank[235] ), .B(n32), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n373 ) );
  MX2X1 U1150 ( .A(\iRF_stage/reg_bank/reg_bank[234] ), .B(n33), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n372 ) );
  MX2X1 U1151 ( .A(\iRF_stage/reg_bank/reg_bank[233] ), .B(n3), .S0(n631), .Y(
        \iRF_stage/reg_bank/n371 ) );
  MX2X1 U1152 ( .A(\iRF_stage/reg_bank/reg_bank[232] ), .B(n4), .S0(n631), .Y(
        \iRF_stage/reg_bank/n370 ) );
  MX2X1 U1153 ( .A(\iRF_stage/reg_bank/reg_bank[231] ), .B(n5), .S0(n631), .Y(
        \iRF_stage/reg_bank/n369 ) );
  MX2X1 U1154 ( .A(\iRF_stage/reg_bank/reg_bank[230] ), .B(n6), .S0(n631), .Y(
        \iRF_stage/reg_bank/n368 ) );
  MX2X1 U1155 ( .A(\iRF_stage/reg_bank/reg_bank[229] ), .B(n7), .S0(n631), .Y(
        \iRF_stage/reg_bank/n367 ) );
  MX2X1 U1156 ( .A(\iRF_stage/reg_bank/reg_bank[228] ), .B(n8), .S0(n631), .Y(
        \iRF_stage/reg_bank/n366 ) );
  MX2X1 U1157 ( .A(\iRF_stage/reg_bank/reg_bank[227] ), .B(n9), .S0(n631), .Y(
        \iRF_stage/reg_bank/n365 ) );
  MX2X1 U1158 ( .A(\iRF_stage/reg_bank/reg_bank[226] ), .B(n12), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n364 ) );
  MX2X1 U1159 ( .A(\iRF_stage/reg_bank/reg_bank[225] ), .B(n23), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n363 ) );
  MX2X1 U1160 ( .A(\iRF_stage/reg_bank/reg_bank[224] ), .B(n34), .S0(n631), 
        .Y(\iRF_stage/reg_bank/n362 ) );
  AND2X1 U1161 ( .A(n632), .B(n606), .Y(n631) );
  MX2X1 U1162 ( .A(\iRF_stage/reg_bank/reg_bank[223] ), .B(n10), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n361 ) );
  MX2X1 U1163 ( .A(\iRF_stage/reg_bank/reg_bank[222] ), .B(n11), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n360 ) );
  MX2X1 U1164 ( .A(\iRF_stage/reg_bank/reg_bank[221] ), .B(n13), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n359 ) );
  MX2X1 U1165 ( .A(\iRF_stage/reg_bank/reg_bank[220] ), .B(n14), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n358 ) );
  MX2X1 U1166 ( .A(\iRF_stage/reg_bank/reg_bank[219] ), .B(n15), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n357 ) );
  MX2X1 U1167 ( .A(\iRF_stage/reg_bank/reg_bank[218] ), .B(n16), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n356 ) );
  MX2X1 U1168 ( .A(\iRF_stage/reg_bank/reg_bank[217] ), .B(n17), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n355 ) );
  MX2X1 U1169 ( .A(\iRF_stage/reg_bank/reg_bank[216] ), .B(n18), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n354 ) );
  MX2X1 U1170 ( .A(\iRF_stage/reg_bank/reg_bank[215] ), .B(n19), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n353 ) );
  MX2X1 U1171 ( .A(\iRF_stage/reg_bank/reg_bank[214] ), .B(n20), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n352 ) );
  MX2X1 U1172 ( .A(\iRF_stage/reg_bank/reg_bank[213] ), .B(n21), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n351 ) );
  MX2X1 U1173 ( .A(\iRF_stage/reg_bank/reg_bank[212] ), .B(n22), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n350 ) );
  MX2X1 U1174 ( .A(\iRF_stage/reg_bank/reg_bank[211] ), .B(n24), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n349 ) );
  MX2X1 U1175 ( .A(\iRF_stage/reg_bank/reg_bank[210] ), .B(n25), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n348 ) );
  MX2X1 U1176 ( .A(\iRF_stage/reg_bank/reg_bank[209] ), .B(n26), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n347 ) );
  MX2X1 U1177 ( .A(\iRF_stage/reg_bank/reg_bank[208] ), .B(n27), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n346 ) );
  MX2X1 U1178 ( .A(\iRF_stage/reg_bank/reg_bank[207] ), .B(n28), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n345 ) );
  MX2X1 U1179 ( .A(\iRF_stage/reg_bank/reg_bank[206] ), .B(n29), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n344 ) );
  MX2X1 U1180 ( .A(\iRF_stage/reg_bank/reg_bank[205] ), .B(n30), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n343 ) );
  MX2X1 U1181 ( .A(\iRF_stage/reg_bank/reg_bank[204] ), .B(n31), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n342 ) );
  MX2X1 U1182 ( .A(\iRF_stage/reg_bank/reg_bank[203] ), .B(n32), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n341 ) );
  MX2X1 U1183 ( .A(\iRF_stage/reg_bank/reg_bank[202] ), .B(n33), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n340 ) );
  MX2X1 U1184 ( .A(\iRF_stage/reg_bank/reg_bank[201] ), .B(n3), .S0(n633), .Y(
        \iRF_stage/reg_bank/n339 ) );
  MX2X1 U1185 ( .A(\iRF_stage/reg_bank/reg_bank[200] ), .B(n4), .S0(n633), .Y(
        \iRF_stage/reg_bank/n338 ) );
  MX2X1 U1186 ( .A(\iRF_stage/reg_bank/reg_bank[199] ), .B(n5), .S0(n633), .Y(
        \iRF_stage/reg_bank/n337 ) );
  MX2X1 U1187 ( .A(\iRF_stage/reg_bank/reg_bank[198] ), .B(n6), .S0(n633), .Y(
        \iRF_stage/reg_bank/n336 ) );
  MX2X1 U1188 ( .A(\iRF_stage/reg_bank/reg_bank[197] ), .B(n7), .S0(n633), .Y(
        \iRF_stage/reg_bank/n335 ) );
  MX2X1 U1189 ( .A(\iRF_stage/reg_bank/reg_bank[196] ), .B(n8), .S0(n633), .Y(
        \iRF_stage/reg_bank/n334 ) );
  MX2X1 U1190 ( .A(\iRF_stage/reg_bank/reg_bank[195] ), .B(n9), .S0(n633), .Y(
        \iRF_stage/reg_bank/n333 ) );
  MX2X1 U1191 ( .A(\iRF_stage/reg_bank/reg_bank[194] ), .B(n12), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n332 ) );
  MX2X1 U1192 ( .A(\iRF_stage/reg_bank/reg_bank[193] ), .B(n23), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n331 ) );
  MX2X1 U1193 ( .A(\iRF_stage/reg_bank/reg_bank[192] ), .B(n34), .S0(n633), 
        .Y(\iRF_stage/reg_bank/n330 ) );
  AND2X1 U1194 ( .A(n632), .B(n609), .Y(n633) );
  MX2X1 U1195 ( .A(\iRF_stage/reg_bank/reg_bank[191] ), .B(n10), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n329 ) );
  MX2X1 U1196 ( .A(\iRF_stage/reg_bank/reg_bank[190] ), .B(n11), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n328 ) );
  MX2X1 U1197 ( .A(\iRF_stage/reg_bank/reg_bank[189] ), .B(n13), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n327 ) );
  MX2X1 U1198 ( .A(\iRF_stage/reg_bank/reg_bank[188] ), .B(n14), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n326 ) );
  MX2X1 U1199 ( .A(\iRF_stage/reg_bank/reg_bank[187] ), .B(n15), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n325 ) );
  MX2X1 U1200 ( .A(\iRF_stage/reg_bank/reg_bank[186] ), .B(n16), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n324 ) );
  MX2X1 U1201 ( .A(\iRF_stage/reg_bank/reg_bank[185] ), .B(n17), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n323 ) );
  MX2X1 U1202 ( .A(\iRF_stage/reg_bank/reg_bank[184] ), .B(n18), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n322 ) );
  MX2X1 U1203 ( .A(\iRF_stage/reg_bank/reg_bank[183] ), .B(n19), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n321 ) );
  MX2X1 U1204 ( .A(\iRF_stage/reg_bank/reg_bank[182] ), .B(n20), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n320 ) );
  MX2X1 U1205 ( .A(\iRF_stage/reg_bank/reg_bank[181] ), .B(n21), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n319 ) );
  MX2X1 U1206 ( .A(\iRF_stage/reg_bank/reg_bank[180] ), .B(n22), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n318 ) );
  MX2X1 U1207 ( .A(\iRF_stage/reg_bank/reg_bank[179] ), .B(n24), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n317 ) );
  MX2X1 U1208 ( .A(\iRF_stage/reg_bank/reg_bank[178] ), .B(n25), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n316 ) );
  MX2X1 U1209 ( .A(\iRF_stage/reg_bank/reg_bank[177] ), .B(n26), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n315 ) );
  MX2X1 U1210 ( .A(\iRF_stage/reg_bank/reg_bank[176] ), .B(n27), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n314 ) );
  MX2X1 U1211 ( .A(\iRF_stage/reg_bank/reg_bank[175] ), .B(n28), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n313 ) );
  MX2X1 U1212 ( .A(\iRF_stage/reg_bank/reg_bank[174] ), .B(n29), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n312 ) );
  MX2X1 U1213 ( .A(\iRF_stage/reg_bank/reg_bank[173] ), .B(n30), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n311 ) );
  MX2X1 U1214 ( .A(\iRF_stage/reg_bank/reg_bank[172] ), .B(n31), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n310 ) );
  MX2X1 U1215 ( .A(\iRF_stage/reg_bank/reg_bank[171] ), .B(n32), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n309 ) );
  MX2X1 U1216 ( .A(\iRF_stage/reg_bank/reg_bank[170] ), .B(n33), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n308 ) );
  MX2X1 U1217 ( .A(\iRF_stage/reg_bank/reg_bank[169] ), .B(n3), .S0(n634), .Y(
        \iRF_stage/reg_bank/n307 ) );
  MX2X1 U1218 ( .A(\iRF_stage/reg_bank/reg_bank[168] ), .B(n4), .S0(n634), .Y(
        \iRF_stage/reg_bank/n306 ) );
  MX2X1 U1219 ( .A(\iRF_stage/reg_bank/reg_bank[167] ), .B(n5), .S0(n634), .Y(
        \iRF_stage/reg_bank/n305 ) );
  MX2X1 U1220 ( .A(\iRF_stage/reg_bank/reg_bank[166] ), .B(n6), .S0(n634), .Y(
        \iRF_stage/reg_bank/n304 ) );
  MX2X1 U1221 ( .A(\iRF_stage/reg_bank/reg_bank[165] ), .B(n7), .S0(n634), .Y(
        \iRF_stage/reg_bank/n303 ) );
  MX2X1 U1222 ( .A(\iRF_stage/reg_bank/reg_bank[164] ), .B(n8), .S0(n634), .Y(
        \iRF_stage/reg_bank/n302 ) );
  MX2X1 U1223 ( .A(\iRF_stage/reg_bank/reg_bank[163] ), .B(n9), .S0(n634), .Y(
        \iRF_stage/reg_bank/n301 ) );
  MX2X1 U1224 ( .A(\iRF_stage/reg_bank/reg_bank[162] ), .B(n12), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n300 ) );
  MX2X1 U1225 ( .A(\iRF_stage/reg_bank/reg_bank[161] ), .B(n23), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n299 ) );
  MX2X1 U1226 ( .A(\iRF_stage/reg_bank/reg_bank[160] ), .B(n34), .S0(n634), 
        .Y(\iRF_stage/reg_bank/n298 ) );
  AND2X1 U1227 ( .A(n632), .B(n611), .Y(n634) );
  MX2X1 U1228 ( .A(\iRF_stage/reg_bank/reg_bank[159] ), .B(n10), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n297 ) );
  MX2X1 U1229 ( .A(\iRF_stage/reg_bank/reg_bank[158] ), .B(n11), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n296 ) );
  MX2X1 U1230 ( .A(\iRF_stage/reg_bank/reg_bank[157] ), .B(n13), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n295 ) );
  MX2X1 U1231 ( .A(\iRF_stage/reg_bank/reg_bank[156] ), .B(n14), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n294 ) );
  MX2X1 U1232 ( .A(\iRF_stage/reg_bank/reg_bank[155] ), .B(n15), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n293 ) );
  MX2X1 U1233 ( .A(\iRF_stage/reg_bank/reg_bank[154] ), .B(n16), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n292 ) );
  MX2X1 U1234 ( .A(\iRF_stage/reg_bank/reg_bank[153] ), .B(n17), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n291 ) );
  MX2X1 U1235 ( .A(\iRF_stage/reg_bank/reg_bank[152] ), .B(n18), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n290 ) );
  MX2X1 U1236 ( .A(\iRF_stage/reg_bank/reg_bank[151] ), .B(n19), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n289 ) );
  MX2X1 U1237 ( .A(\iRF_stage/reg_bank/reg_bank[150] ), .B(n20), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n288 ) );
  MX2X1 U1238 ( .A(\iRF_stage/reg_bank/reg_bank[149] ), .B(n21), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n287 ) );
  MX2X1 U1239 ( .A(\iRF_stage/reg_bank/reg_bank[148] ), .B(n22), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n286 ) );
  MX2X1 U1240 ( .A(\iRF_stage/reg_bank/reg_bank[147] ), .B(n24), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n285 ) );
  MX2X1 U1241 ( .A(\iRF_stage/reg_bank/reg_bank[146] ), .B(n25), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n284 ) );
  MX2X1 U1242 ( .A(\iRF_stage/reg_bank/reg_bank[145] ), .B(n26), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n283 ) );
  MX2X1 U1243 ( .A(\iRF_stage/reg_bank/reg_bank[144] ), .B(n27), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n282 ) );
  MX2X1 U1244 ( .A(\iRF_stage/reg_bank/reg_bank[143] ), .B(n28), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n281 ) );
  MX2X1 U1245 ( .A(\iRF_stage/reg_bank/reg_bank[142] ), .B(n29), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n280 ) );
  MX2X1 U1246 ( .A(\iRF_stage/reg_bank/reg_bank[141] ), .B(n30), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n279 ) );
  MX2X1 U1247 ( .A(\iRF_stage/reg_bank/reg_bank[140] ), .B(n31), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n278 ) );
  MX2X1 U1248 ( .A(\iRF_stage/reg_bank/reg_bank[139] ), .B(n32), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n277 ) );
  MX2X1 U1249 ( .A(\iRF_stage/reg_bank/reg_bank[138] ), .B(n33), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n276 ) );
  MX2X1 U1250 ( .A(\iRF_stage/reg_bank/reg_bank[137] ), .B(n3), .S0(n635), .Y(
        \iRF_stage/reg_bank/n275 ) );
  MX2X1 U1251 ( .A(\iRF_stage/reg_bank/reg_bank[136] ), .B(n4), .S0(n635), .Y(
        \iRF_stage/reg_bank/n274 ) );
  MX2X1 U1252 ( .A(\iRF_stage/reg_bank/reg_bank[135] ), .B(n5), .S0(n635), .Y(
        \iRF_stage/reg_bank/n273 ) );
  MX2X1 U1253 ( .A(\iRF_stage/reg_bank/reg_bank[134] ), .B(n6), .S0(n635), .Y(
        \iRF_stage/reg_bank/n272 ) );
  MX2X1 U1254 ( .A(\iRF_stage/reg_bank/reg_bank[133] ), .B(n7), .S0(n635), .Y(
        \iRF_stage/reg_bank/n271 ) );
  MX2X1 U1255 ( .A(\iRF_stage/reg_bank/reg_bank[132] ), .B(n8), .S0(n635), .Y(
        \iRF_stage/reg_bank/n270 ) );
  MX2X1 U1256 ( .A(\iRF_stage/reg_bank/reg_bank[131] ), .B(n9), .S0(n635), .Y(
        \iRF_stage/reg_bank/n269 ) );
  MX2X1 U1257 ( .A(\iRF_stage/reg_bank/reg_bank[130] ), .B(n12), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n268 ) );
  MX2X1 U1258 ( .A(\iRF_stage/reg_bank/reg_bank[129] ), .B(n23), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n267 ) );
  MX2X1 U1259 ( .A(\iRF_stage/reg_bank/reg_bank[128] ), .B(n34), .S0(n635), 
        .Y(\iRF_stage/reg_bank/n266 ) );
  AND2X1 U1260 ( .A(n632), .B(n613), .Y(n635) );
  MX2X1 U1261 ( .A(\iRF_stage/reg_bank/reg_bank[127] ), .B(n10), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n265 ) );
  MX2X1 U1262 ( .A(\iRF_stage/reg_bank/reg_bank[126] ), .B(n11), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n264 ) );
  MX2X1 U1263 ( .A(\iRF_stage/reg_bank/reg_bank[125] ), .B(n13), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n263 ) );
  MX2X1 U1264 ( .A(\iRF_stage/reg_bank/reg_bank[124] ), .B(n14), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n262 ) );
  MX2X1 U1265 ( .A(\iRF_stage/reg_bank/reg_bank[123] ), .B(n15), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n261 ) );
  MX2X1 U1266 ( .A(\iRF_stage/reg_bank/reg_bank[122] ), .B(n16), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n260 ) );
  MX2X1 U1267 ( .A(\iRF_stage/reg_bank/reg_bank[121] ), .B(n17), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n259 ) );
  MX2X1 U1268 ( .A(\iRF_stage/reg_bank/reg_bank[120] ), .B(n18), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n258 ) );
  MX2X1 U1269 ( .A(\iRF_stage/reg_bank/reg_bank[119] ), .B(n19), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n257 ) );
  MX2X1 U1270 ( .A(\iRF_stage/reg_bank/reg_bank[118] ), .B(n20), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n256 ) );
  MX2X1 U1271 ( .A(\iRF_stage/reg_bank/reg_bank[117] ), .B(n21), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n255 ) );
  MX2X1 U1272 ( .A(\iRF_stage/reg_bank/reg_bank[116] ), .B(n22), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n254 ) );
  MX2X1 U1273 ( .A(\iRF_stage/reg_bank/reg_bank[115] ), .B(n24), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n253 ) );
  MX2X1 U1274 ( .A(\iRF_stage/reg_bank/reg_bank[114] ), .B(n25), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n252 ) );
  MX2X1 U1275 ( .A(\iRF_stage/reg_bank/reg_bank[113] ), .B(n26), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n251 ) );
  MX2X1 U1276 ( .A(\iRF_stage/reg_bank/reg_bank[112] ), .B(n27), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n250 ) );
  MX2X1 U1277 ( .A(\iRF_stage/reg_bank/reg_bank[111] ), .B(n28), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n249 ) );
  MX2X1 U1278 ( .A(\iRF_stage/reg_bank/reg_bank[110] ), .B(n29), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n248 ) );
  MX2X1 U1279 ( .A(\iRF_stage/reg_bank/reg_bank[109] ), .B(n30), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n247 ) );
  MX2X1 U1280 ( .A(\iRF_stage/reg_bank/reg_bank[108] ), .B(n31), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n246 ) );
  MX2X1 U1281 ( .A(\iRF_stage/reg_bank/reg_bank[107] ), .B(n32), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n245 ) );
  MX2X1 U1282 ( .A(\iRF_stage/reg_bank/reg_bank[106] ), .B(n33), .S0(n636), 
        .Y(\iRF_stage/reg_bank/n244 ) );
  MX2X1 U1283 ( .A(\iRF_stage/reg_bank/reg_bank[105] ), .B(n3), .S0(n636), .Y(
        \iRF_stage/reg_bank/n243 ) );
  MX2X1 U1284 ( .A(\iRF_stage/reg_bank/reg_bank[104] ), .B(n4), .S0(n636), .Y(
        \iRF_stage/reg_bank/n242 ) );
  MX2X1 U1285 ( .A(\iRF_stage/reg_bank/reg_bank[103] ), .B(n5), .S0(n636), .Y(
        \iRF_stage/reg_bank/n241 ) );
  MX2X1 U1286 ( .A(\iRF_stage/reg_bank/reg_bank[102] ), .B(n6), .S0(n636), .Y(
        \iRF_stage/reg_bank/n240 ) );
  MX2X1 U1287 ( .A(\iRF_stage/reg_bank/reg_bank[101] ), .B(n7), .S0(n636), .Y(
        \iRF_stage/reg_bank/n239 ) );
  MX2X1 U1288 ( .A(\iRF_stage/reg_bank/reg_bank[100] ), .B(n8), .S0(n636), .Y(
        \iRF_stage/reg_bank/n238 ) );
  MX2X1 U1289 ( .A(\iRF_stage/reg_bank/reg_bank[99] ), .B(n9), .S0(n636), .Y(
        \iRF_stage/reg_bank/n237 ) );
  MX2X1 U1290 ( .A(\iRF_stage/reg_bank/reg_bank[98] ), .B(n12), .S0(n636), .Y(
        \iRF_stage/reg_bank/n236 ) );
  MX2X1 U1291 ( .A(\iRF_stage/reg_bank/reg_bank[97] ), .B(n23), .S0(n636), .Y(
        \iRF_stage/reg_bank/n235 ) );
  MX2X1 U1292 ( .A(\iRF_stage/reg_bank/reg_bank[96] ), .B(n34), .S0(n636), .Y(
        \iRF_stage/reg_bank/n234 ) );
  AND2X1 U1293 ( .A(n632), .B(n615), .Y(n636) );
  MX2X1 U1294 ( .A(\iRF_stage/reg_bank/reg_bank[95] ), .B(n10), .S0(n637), .Y(
        \iRF_stage/reg_bank/n233 ) );
  MX2X1 U1295 ( .A(\iRF_stage/reg_bank/reg_bank[94] ), .B(n11), .S0(n637), .Y(
        \iRF_stage/reg_bank/n232 ) );
  MX2X1 U1296 ( .A(\iRF_stage/reg_bank/reg_bank[93] ), .B(n13), .S0(n637), .Y(
        \iRF_stage/reg_bank/n231 ) );
  MX2X1 U1297 ( .A(\iRF_stage/reg_bank/reg_bank[92] ), .B(n14), .S0(n637), .Y(
        \iRF_stage/reg_bank/n230 ) );
  MX2X1 U1298 ( .A(\iRF_stage/reg_bank/reg_bank[91] ), .B(n15), .S0(n637), .Y(
        \iRF_stage/reg_bank/n229 ) );
  MX2X1 U1299 ( .A(\iRF_stage/reg_bank/reg_bank[90] ), .B(n16), .S0(n637), .Y(
        \iRF_stage/reg_bank/n228 ) );
  MX2X1 U1300 ( .A(\iRF_stage/reg_bank/reg_bank[89] ), .B(n17), .S0(n637), .Y(
        \iRF_stage/reg_bank/n227 ) );
  MX2X1 U1301 ( .A(\iRF_stage/reg_bank/reg_bank[88] ), .B(n18), .S0(n637), .Y(
        \iRF_stage/reg_bank/n226 ) );
  MX2X1 U1302 ( .A(\iRF_stage/reg_bank/reg_bank[87] ), .B(n19), .S0(n637), .Y(
        \iRF_stage/reg_bank/n225 ) );
  MX2X1 U1303 ( .A(\iRF_stage/reg_bank/reg_bank[86] ), .B(n20), .S0(n637), .Y(
        \iRF_stage/reg_bank/n224 ) );
  MX2X1 U1304 ( .A(\iRF_stage/reg_bank/reg_bank[85] ), .B(n21), .S0(n637), .Y(
        \iRF_stage/reg_bank/n223 ) );
  MX2X1 U1305 ( .A(\iRF_stage/reg_bank/reg_bank[84] ), .B(n22), .S0(n637), .Y(
        \iRF_stage/reg_bank/n222 ) );
  MX2X1 U1306 ( .A(\iRF_stage/reg_bank/reg_bank[83] ), .B(n24), .S0(n637), .Y(
        \iRF_stage/reg_bank/n221 ) );
  MX2X1 U1307 ( .A(\iRF_stage/reg_bank/reg_bank[82] ), .B(n25), .S0(n637), .Y(
        \iRF_stage/reg_bank/n220 ) );
  MX2X1 U1308 ( .A(\iRF_stage/reg_bank/reg_bank[81] ), .B(n26), .S0(n637), .Y(
        \iRF_stage/reg_bank/n219 ) );
  MX2X1 U1309 ( .A(\iRF_stage/reg_bank/reg_bank[80] ), .B(n27), .S0(n637), .Y(
        \iRF_stage/reg_bank/n218 ) );
  MX2X1 U1310 ( .A(\iRF_stage/reg_bank/reg_bank[79] ), .B(n28), .S0(n637), .Y(
        \iRF_stage/reg_bank/n217 ) );
  MX2X1 U1311 ( .A(\iRF_stage/reg_bank/reg_bank[78] ), .B(n29), .S0(n637), .Y(
        \iRF_stage/reg_bank/n216 ) );
  MX2X1 U1312 ( .A(\iRF_stage/reg_bank/reg_bank[77] ), .B(n30), .S0(n637), .Y(
        \iRF_stage/reg_bank/n215 ) );
  MX2X1 U1313 ( .A(\iRF_stage/reg_bank/reg_bank[76] ), .B(n31), .S0(n637), .Y(
        \iRF_stage/reg_bank/n214 ) );
  MX2X1 U1314 ( .A(\iRF_stage/reg_bank/reg_bank[75] ), .B(n32), .S0(n637), .Y(
        \iRF_stage/reg_bank/n213 ) );
  MX2X1 U1315 ( .A(\iRF_stage/reg_bank/reg_bank[74] ), .B(n33), .S0(n637), .Y(
        \iRF_stage/reg_bank/n212 ) );
  MX2X1 U1316 ( .A(\iRF_stage/reg_bank/reg_bank[73] ), .B(n3), .S0(n637), .Y(
        \iRF_stage/reg_bank/n211 ) );
  MX2X1 U1317 ( .A(\iRF_stage/reg_bank/reg_bank[72] ), .B(n4), .S0(n637), .Y(
        \iRF_stage/reg_bank/n210 ) );
  MX2X1 U1318 ( .A(\iRF_stage/reg_bank/reg_bank[71] ), .B(n5), .S0(n637), .Y(
        \iRF_stage/reg_bank/n209 ) );
  MX2X1 U1319 ( .A(\iRF_stage/reg_bank/reg_bank[70] ), .B(n6), .S0(n637), .Y(
        \iRF_stage/reg_bank/n208 ) );
  MX2X1 U1320 ( .A(\iRF_stage/reg_bank/reg_bank[69] ), .B(n7), .S0(n637), .Y(
        \iRF_stage/reg_bank/n207 ) );
  MX2X1 U1321 ( .A(\iRF_stage/reg_bank/reg_bank[68] ), .B(n8), .S0(n637), .Y(
        \iRF_stage/reg_bank/n206 ) );
  MX2X1 U1322 ( .A(\iRF_stage/reg_bank/reg_bank[67] ), .B(n9), .S0(n637), .Y(
        \iRF_stage/reg_bank/n205 ) );
  MX2X1 U1323 ( .A(\iRF_stage/reg_bank/reg_bank[66] ), .B(n12), .S0(n637), .Y(
        \iRF_stage/reg_bank/n204 ) );
  MX2X1 U1324 ( .A(\iRF_stage/reg_bank/reg_bank[65] ), .B(n23), .S0(n637), .Y(
        \iRF_stage/reg_bank/n203 ) );
  MX2X1 U1325 ( .A(\iRF_stage/reg_bank/reg_bank[64] ), .B(n34), .S0(n637), .Y(
        \iRF_stage/reg_bank/n202 ) );
  AND2X1 U1326 ( .A(n632), .B(n617), .Y(n637) );
  MX2X1 U1327 ( .A(\iRF_stage/reg_bank/reg_bank[63] ), .B(n10), .S0(n638), .Y(
        \iRF_stage/reg_bank/n201 ) );
  MX2X1 U1328 ( .A(\iRF_stage/reg_bank/reg_bank[62] ), .B(n11), .S0(n638), .Y(
        \iRF_stage/reg_bank/n200 ) );
  MX2X1 U1329 ( .A(\iRF_stage/reg_bank/reg_bank[61] ), .B(n13), .S0(n638), .Y(
        \iRF_stage/reg_bank/n199 ) );
  MX2X1 U1330 ( .A(\iRF_stage/reg_bank/reg_bank[60] ), .B(n14), .S0(n638), .Y(
        \iRF_stage/reg_bank/n198 ) );
  MX2X1 U1331 ( .A(\iRF_stage/reg_bank/reg_bank[59] ), .B(n15), .S0(n638), .Y(
        \iRF_stage/reg_bank/n197 ) );
  MX2X1 U1332 ( .A(\iRF_stage/reg_bank/reg_bank[58] ), .B(n16), .S0(n638), .Y(
        \iRF_stage/reg_bank/n196 ) );
  MX2X1 U1333 ( .A(\iRF_stage/reg_bank/reg_bank[57] ), .B(n17), .S0(n638), .Y(
        \iRF_stage/reg_bank/n195 ) );
  MX2X1 U1334 ( .A(\iRF_stage/reg_bank/reg_bank[56] ), .B(n18), .S0(n638), .Y(
        \iRF_stage/reg_bank/n194 ) );
  MX2X1 U1335 ( .A(\iRF_stage/reg_bank/reg_bank[55] ), .B(n19), .S0(n638), .Y(
        \iRF_stage/reg_bank/n193 ) );
  MX2X1 U1336 ( .A(\iRF_stage/reg_bank/reg_bank[54] ), .B(n20), .S0(n638), .Y(
        \iRF_stage/reg_bank/n192 ) );
  MX2X1 U1337 ( .A(\iRF_stage/reg_bank/reg_bank[53] ), .B(n21), .S0(n638), .Y(
        \iRF_stage/reg_bank/n191 ) );
  MX2X1 U1338 ( .A(\iRF_stage/reg_bank/reg_bank[52] ), .B(n22), .S0(n638), .Y(
        \iRF_stage/reg_bank/n190 ) );
  MX2X1 U1339 ( .A(\iRF_stage/reg_bank/reg_bank[51] ), .B(n24), .S0(n638), .Y(
        \iRF_stage/reg_bank/n189 ) );
  MX2X1 U1340 ( .A(\iRF_stage/reg_bank/reg_bank[50] ), .B(n25), .S0(n638), .Y(
        \iRF_stage/reg_bank/n188 ) );
  MX2X1 U1341 ( .A(\iRF_stage/reg_bank/reg_bank[49] ), .B(n26), .S0(n638), .Y(
        \iRF_stage/reg_bank/n187 ) );
  MX2X1 U1342 ( .A(\iRF_stage/reg_bank/reg_bank[48] ), .B(n27), .S0(n638), .Y(
        \iRF_stage/reg_bank/n186 ) );
  MX2X1 U1343 ( .A(\iRF_stage/reg_bank/reg_bank[47] ), .B(n28), .S0(n638), .Y(
        \iRF_stage/reg_bank/n185 ) );
  MX2X1 U1344 ( .A(\iRF_stage/reg_bank/reg_bank[46] ), .B(n29), .S0(n638), .Y(
        \iRF_stage/reg_bank/n184 ) );
  MX2X1 U1345 ( .A(\iRF_stage/reg_bank/reg_bank[45] ), .B(n30), .S0(n638), .Y(
        \iRF_stage/reg_bank/n183 ) );
  MX2X1 U1346 ( .A(\iRF_stage/reg_bank/reg_bank[44] ), .B(n31), .S0(n638), .Y(
        \iRF_stage/reg_bank/n182 ) );
  MX2X1 U1347 ( .A(\iRF_stage/reg_bank/reg_bank[43] ), .B(n32), .S0(n638), .Y(
        \iRF_stage/reg_bank/n181 ) );
  MX2X1 U1348 ( .A(\iRF_stage/reg_bank/reg_bank[42] ), .B(n33), .S0(n638), .Y(
        \iRF_stage/reg_bank/n180 ) );
  MX2X1 U1349 ( .A(\iRF_stage/reg_bank/reg_bank[41] ), .B(n3), .S0(n638), .Y(
        \iRF_stage/reg_bank/n179 ) );
  MX2X1 U1350 ( .A(\iRF_stage/reg_bank/reg_bank[40] ), .B(n4), .S0(n638), .Y(
        \iRF_stage/reg_bank/n178 ) );
  MX2X1 U1351 ( .A(\iRF_stage/reg_bank/reg_bank[39] ), .B(n5), .S0(n638), .Y(
        \iRF_stage/reg_bank/n177 ) );
  MX2X1 U1352 ( .A(\iRF_stage/reg_bank/reg_bank[38] ), .B(n6), .S0(n638), .Y(
        \iRF_stage/reg_bank/n176 ) );
  MX2X1 U1353 ( .A(\iRF_stage/reg_bank/reg_bank[37] ), .B(n7), .S0(n638), .Y(
        \iRF_stage/reg_bank/n175 ) );
  MX2X1 U1354 ( .A(\iRF_stage/reg_bank/reg_bank[36] ), .B(n8), .S0(n638), .Y(
        \iRF_stage/reg_bank/n174 ) );
  MX2X1 U1355 ( .A(\iRF_stage/reg_bank/reg_bank[35] ), .B(n9), .S0(n638), .Y(
        \iRF_stage/reg_bank/n173 ) );
  MX2X1 U1356 ( .A(\iRF_stage/reg_bank/reg_bank[34] ), .B(n12), .S0(n638), .Y(
        \iRF_stage/reg_bank/n172 ) );
  MX2X1 U1357 ( .A(\iRF_stage/reg_bank/reg_bank[33] ), .B(n23), .S0(n638), .Y(
        \iRF_stage/reg_bank/n171 ) );
  MX2X1 U1358 ( .A(\iRF_stage/reg_bank/reg_bank[32] ), .B(n34), .S0(n638), .Y(
        \iRF_stage/reg_bank/n170 ) );
  AND2X1 U1359 ( .A(n632), .B(n601), .Y(n638) );
  NOR3X1 U1360 ( .A(n639), .B(\iRF_stage/reg_bank/r_wraddress[0] ), .C(n640), 
        .Y(n601) );
  MX2X1 U1361 ( .A(\iRF_stage/reg_bank/reg_bank[31] ), .B(n10), .S0(n641), .Y(
        \iRF_stage/reg_bank/n169 ) );
  MX2X1 U1362 ( .A(\iRF_stage/reg_bank/reg_bank[30] ), .B(n11), .S0(n641), .Y(
        \iRF_stage/reg_bank/n168 ) );
  MX2X1 U1363 ( .A(\iRF_stage/reg_bank/reg_bank[29] ), .B(n13), .S0(n641), .Y(
        \iRF_stage/reg_bank/n167 ) );
  MX2X1 U1364 ( .A(\iRF_stage/reg_bank/reg_bank[28] ), .B(n14), .S0(n641), .Y(
        \iRF_stage/reg_bank/n166 ) );
  MX2X1 U1365 ( .A(\iRF_stage/reg_bank/reg_bank[27] ), .B(n15), .S0(n641), .Y(
        \iRF_stage/reg_bank/n165 ) );
  MX2X1 U1366 ( .A(\iRF_stage/reg_bank/reg_bank[26] ), .B(n16), .S0(n641), .Y(
        \iRF_stage/reg_bank/n164 ) );
  MX2X1 U1367 ( .A(\iRF_stage/reg_bank/reg_bank[25] ), .B(n17), .S0(n641), .Y(
        \iRF_stage/reg_bank/n163 ) );
  MX2X1 U1368 ( .A(\iRF_stage/reg_bank/reg_bank[24] ), .B(n18), .S0(n641), .Y(
        \iRF_stage/reg_bank/n162 ) );
  MX2X1 U1369 ( .A(\iRF_stage/reg_bank/reg_bank[23] ), .B(n19), .S0(n641), .Y(
        \iRF_stage/reg_bank/n161 ) );
  MX2X1 U1370 ( .A(\iRF_stage/reg_bank/reg_bank[22] ), .B(n20), .S0(n641), .Y(
        \iRF_stage/reg_bank/n160 ) );
  MX2X1 U1371 ( .A(\iRF_stage/reg_bank/reg_bank[21] ), .B(n21), .S0(n641), .Y(
        \iRF_stage/reg_bank/n159 ) );
  MX2X1 U1372 ( .A(\iRF_stage/reg_bank/reg_bank[20] ), .B(n22), .S0(n641), .Y(
        \iRF_stage/reg_bank/n158 ) );
  MX2X1 U1373 ( .A(\iRF_stage/reg_bank/reg_bank[19] ), .B(n24), .S0(n641), .Y(
        \iRF_stage/reg_bank/n157 ) );
  MX2X1 U1374 ( .A(\iRF_stage/reg_bank/reg_bank[18] ), .B(n25), .S0(n641), .Y(
        \iRF_stage/reg_bank/n156 ) );
  MX2X1 U1375 ( .A(\iRF_stage/reg_bank/reg_bank[17] ), .B(n26), .S0(n641), .Y(
        \iRF_stage/reg_bank/n155 ) );
  MX2X1 U1376 ( .A(\iRF_stage/reg_bank/reg_bank[16] ), .B(n27), .S0(n641), .Y(
        \iRF_stage/reg_bank/n154 ) );
  MX2X1 U1377 ( .A(\iRF_stage/reg_bank/reg_bank[15] ), .B(n28), .S0(n641), .Y(
        \iRF_stage/reg_bank/n153 ) );
  MX2X1 U1378 ( .A(\iRF_stage/reg_bank/reg_bank[14] ), .B(n29), .S0(n641), .Y(
        \iRF_stage/reg_bank/n152 ) );
  MX2X1 U1379 ( .A(\iRF_stage/reg_bank/reg_bank[13] ), .B(n30), .S0(n641), .Y(
        \iRF_stage/reg_bank/n151 ) );
  MX2X1 U1380 ( .A(\iRF_stage/reg_bank/reg_bank[12] ), .B(n31), .S0(n641), .Y(
        \iRF_stage/reg_bank/n150 ) );
  MX2X1 U1381 ( .A(\iRF_stage/reg_bank/reg_bank[11] ), .B(n32), .S0(n641), .Y(
        \iRF_stage/reg_bank/n149 ) );
  MX2X1 U1382 ( .A(\iRF_stage/reg_bank/reg_bank[10] ), .B(n33), .S0(n641), .Y(
        \iRF_stage/reg_bank/n148 ) );
  MX2X1 U1383 ( .A(\iRF_stage/reg_bank/reg_bank[9] ), .B(n3), .S0(n641), .Y(
        \iRF_stage/reg_bank/n147 ) );
  MX2X1 U1384 ( .A(\iRF_stage/reg_bank/reg_bank[8] ), .B(n4), .S0(n641), .Y(
        \iRF_stage/reg_bank/n146 ) );
  MX2X1 U1385 ( .A(\iRF_stage/reg_bank/reg_bank[7] ), .B(n5), .S0(n641), .Y(
        \iRF_stage/reg_bank/n145 ) );
  MX2X1 U1386 ( .A(\iRF_stage/reg_bank/reg_bank[6] ), .B(n6), .S0(n641), .Y(
        \iRF_stage/reg_bank/n144 ) );
  MX2X1 U1387 ( .A(\iRF_stage/reg_bank/reg_bank[5] ), .B(n7), .S0(n641), .Y(
        \iRF_stage/reg_bank/n143 ) );
  MX2X1 U1388 ( .A(\iRF_stage/reg_bank/reg_bank[4] ), .B(n8), .S0(n641), .Y(
        \iRF_stage/reg_bank/n142 ) );
  MX2X1 U1389 ( .A(\iRF_stage/reg_bank/reg_bank[3] ), .B(n9), .S0(n641), .Y(
        \iRF_stage/reg_bank/n141 ) );
  MX2X1 U1390 ( .A(\iRF_stage/reg_bank/reg_bank[2] ), .B(n12), .S0(n641), .Y(
        \iRF_stage/reg_bank/n140 ) );
  MX2X1 U1391 ( .A(\iRF_stage/reg_bank/reg_bank[1] ), .B(n23), .S0(n641), .Y(
        \iRF_stage/reg_bank/n139 ) );
  MX2X1 U1392 ( .A(\iRF_stage/reg_bank/reg_bank[0] ), .B(n34), .S0(n641), .Y(
        \iRF_stage/reg_bank/n138 ) );
  AND2X1 U1393 ( .A(n632), .B(n604), .Y(n641) );
  NOR3X1 U1394 ( .A(n642), .B(n639), .C(n640), .Y(n604) );
  NOR3BX1 U1395 ( .AN(\iRF_stage/reg_bank/r_wren ), .B(n620), .C(n630), .Y(
        n632) );
  MX2X1 U1396 ( .A(\iRF_stage/reg_bank/reg_bank[1023] ), .B(n10), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1161 ) );
  MX2X1 U1397 ( .A(\iRF_stage/reg_bank/reg_bank[1022] ), .B(n11), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1160 ) );
  MX2X1 U1398 ( .A(\iRF_stage/reg_bank/reg_bank[1021] ), .B(n13), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1159 ) );
  MX2X1 U1399 ( .A(\iRF_stage/reg_bank/reg_bank[1020] ), .B(n14), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1158 ) );
  MX2X1 U1400 ( .A(\iRF_stage/reg_bank/reg_bank[1019] ), .B(n15), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1157 ) );
  MX2X1 U1401 ( .A(\iRF_stage/reg_bank/reg_bank[1018] ), .B(n16), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1156 ) );
  MX2X1 U1402 ( .A(\iRF_stage/reg_bank/reg_bank[1017] ), .B(n17), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1155 ) );
  MX2X1 U1403 ( .A(\iRF_stage/reg_bank/reg_bank[1016] ), .B(n18), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1154 ) );
  MX2X1 U1404 ( .A(\iRF_stage/reg_bank/reg_bank[1015] ), .B(n19), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1153 ) );
  MX2X1 U1405 ( .A(\iRF_stage/reg_bank/reg_bank[1014] ), .B(n20), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1152 ) );
  MX2X1 U1406 ( .A(\iRF_stage/reg_bank/reg_bank[1013] ), .B(n21), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1151 ) );
  MX2X1 U1407 ( .A(\iRF_stage/reg_bank/reg_bank[1012] ), .B(n22), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1150 ) );
  MX2X1 U1408 ( .A(\iRF_stage/reg_bank/reg_bank[1011] ), .B(n24), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1149 ) );
  MX2X1 U1409 ( .A(\iRF_stage/reg_bank/reg_bank[1010] ), .B(n25), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1148 ) );
  MX2X1 U1410 ( .A(\iRF_stage/reg_bank/reg_bank[1009] ), .B(n26), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1147 ) );
  MX2X1 U1411 ( .A(\iRF_stage/reg_bank/reg_bank[1008] ), .B(n27), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1146 ) );
  MX2X1 U1412 ( .A(\iRF_stage/reg_bank/reg_bank[1007] ), .B(n28), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1145 ) );
  MX2X1 U1413 ( .A(\iRF_stage/reg_bank/reg_bank[1006] ), .B(n29), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1144 ) );
  MX2X1 U1414 ( .A(\iRF_stage/reg_bank/reg_bank[1005] ), .B(n30), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1143 ) );
  MX2X1 U1415 ( .A(\iRF_stage/reg_bank/reg_bank[1004] ), .B(n31), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1142 ) );
  MX2X1 U1416 ( .A(\iRF_stage/reg_bank/reg_bank[1003] ), .B(n32), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1141 ) );
  MX2X1 U1417 ( .A(\iRF_stage/reg_bank/reg_bank[1002] ), .B(n33), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1140 ) );
  MX2X1 U1418 ( .A(\iRF_stage/reg_bank/reg_bank[1001] ), .B(n3), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1139 ) );
  MX2X1 U1419 ( .A(\iRF_stage/reg_bank/reg_bank[1000] ), .B(n4), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1138 ) );
  MX2X1 U1420 ( .A(\iRF_stage/reg_bank/reg_bank[999] ), .B(n5), .S0(n643), .Y(
        \iRF_stage/reg_bank/n1137 ) );
  MX2X1 U1421 ( .A(\iRF_stage/reg_bank/reg_bank[998] ), .B(n6), .S0(n643), .Y(
        \iRF_stage/reg_bank/n1136 ) );
  MX2X1 U1422 ( .A(\iRF_stage/reg_bank/reg_bank[997] ), .B(n7), .S0(n643), .Y(
        \iRF_stage/reg_bank/n1135 ) );
  MX2X1 U1423 ( .A(\iRF_stage/reg_bank/reg_bank[996] ), .B(n8), .S0(n643), .Y(
        \iRF_stage/reg_bank/n1134 ) );
  MX2X1 U1424 ( .A(\iRF_stage/reg_bank/reg_bank[995] ), .B(n9), .S0(n643), .Y(
        \iRF_stage/reg_bank/n1133 ) );
  MX2X1 U1425 ( .A(\iRF_stage/reg_bank/reg_bank[994] ), .B(n12), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1132 ) );
  MX2X1 U1426 ( .A(\iRF_stage/reg_bank/reg_bank[993] ), .B(n23), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1131 ) );
  MX2X1 U1427 ( .A(\iRF_stage/reg_bank/reg_bank[992] ), .B(n34), .S0(n643), 
        .Y(\iRF_stage/reg_bank/n1130 ) );
  AND2X1 U1428 ( .A(n606), .B(n602), .Y(n643) );
  NOR3X1 U1429 ( .A(\iRF_stage/reg_bank/r_wraddress[1] ), .B(
        \iRF_stage/reg_bank/r_wraddress[2] ), .C(
        \iRF_stage/reg_bank/r_wraddress[0] ), .Y(n606) );
  MX2X1 U1430 ( .A(\iRF_stage/reg_bank/reg_bank[991] ), .B(n10), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1129 ) );
  MX2X1 U1431 ( .A(\iRF_stage/reg_bank/reg_bank[990] ), .B(n11), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1128 ) );
  MX2X1 U1432 ( .A(\iRF_stage/reg_bank/reg_bank[989] ), .B(n13), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1127 ) );
  MX2X1 U1433 ( .A(\iRF_stage/reg_bank/reg_bank[988] ), .B(n14), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1126 ) );
  MX2X1 U1434 ( .A(\iRF_stage/reg_bank/reg_bank[987] ), .B(n15), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1125 ) );
  MX2X1 U1435 ( .A(\iRF_stage/reg_bank/reg_bank[986] ), .B(n16), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1124 ) );
  MX2X1 U1436 ( .A(\iRF_stage/reg_bank/reg_bank[985] ), .B(n17), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1123 ) );
  MX2X1 U1437 ( .A(\iRF_stage/reg_bank/reg_bank[984] ), .B(n18), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1122 ) );
  MX2X1 U1438 ( .A(\iRF_stage/reg_bank/reg_bank[983] ), .B(n19), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1121 ) );
  MX2X1 U1439 ( .A(\iRF_stage/reg_bank/reg_bank[982] ), .B(n20), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1120 ) );
  MX2X1 U1440 ( .A(\iRF_stage/reg_bank/reg_bank[981] ), .B(n21), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1119 ) );
  MX2X1 U1441 ( .A(\iRF_stage/reg_bank/reg_bank[980] ), .B(n22), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1118 ) );
  MX2X1 U1442 ( .A(\iRF_stage/reg_bank/reg_bank[979] ), .B(n24), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1117 ) );
  MX2X1 U1443 ( .A(\iRF_stage/reg_bank/reg_bank[978] ), .B(n25), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1116 ) );
  MX2X1 U1444 ( .A(\iRF_stage/reg_bank/reg_bank[977] ), .B(n26), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1115 ) );
  MX2X1 U1445 ( .A(\iRF_stage/reg_bank/reg_bank[976] ), .B(n27), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1114 ) );
  MX2X1 U1446 ( .A(\iRF_stage/reg_bank/reg_bank[975] ), .B(n28), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1113 ) );
  MX2X1 U1447 ( .A(\iRF_stage/reg_bank/reg_bank[974] ), .B(n29), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1112 ) );
  MX2X1 U1448 ( .A(\iRF_stage/reg_bank/reg_bank[973] ), .B(n30), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1111 ) );
  MX2X1 U1449 ( .A(\iRF_stage/reg_bank/reg_bank[972] ), .B(n31), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1110 ) );
  MX2X1 U1450 ( .A(\iRF_stage/reg_bank/reg_bank[971] ), .B(n32), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1109 ) );
  MX2X1 U1451 ( .A(\iRF_stage/reg_bank/reg_bank[970] ), .B(n33), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1108 ) );
  MX2X1 U1452 ( .A(\iRF_stage/reg_bank/reg_bank[969] ), .B(n3), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1107 ) );
  MX2X1 U1453 ( .A(\iRF_stage/reg_bank/reg_bank[968] ), .B(n4), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1106 ) );
  MX2X1 U1454 ( .A(\iRF_stage/reg_bank/reg_bank[967] ), .B(n5), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1105 ) );
  MX2X1 U1455 ( .A(\iRF_stage/reg_bank/reg_bank[966] ), .B(n6), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1104 ) );
  MX2X1 U1456 ( .A(\iRF_stage/reg_bank/reg_bank[965] ), .B(n7), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1103 ) );
  MX2X1 U1457 ( .A(\iRF_stage/reg_bank/reg_bank[964] ), .B(n8), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1102 ) );
  MX2X1 U1458 ( .A(\iRF_stage/reg_bank/reg_bank[963] ), .B(n9), .S0(n644), .Y(
        \iRF_stage/reg_bank/n1101 ) );
  MX2X1 U1459 ( .A(\iRF_stage/reg_bank/reg_bank[962] ), .B(n12), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1100 ) );
  MX2X1 U1460 ( .A(\iRF_stage/reg_bank/reg_bank[961] ), .B(n23), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1099 ) );
  MX2X1 U1461 ( .A(\iRF_stage/reg_bank/reg_bank[960] ), .B(n34), .S0(n644), 
        .Y(\iRF_stage/reg_bank/n1098 ) );
  AND2X1 U1462 ( .A(n609), .B(n602), .Y(n644) );
  NOR3X1 U1463 ( .A(\iRF_stage/reg_bank/r_wraddress[1] ), .B(
        \iRF_stage/reg_bank/r_wraddress[2] ), .C(n642), .Y(n609) );
  MX2X1 U1464 ( .A(\iRF_stage/reg_bank/reg_bank[959] ), .B(n10), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1097 ) );
  MX2X1 U1465 ( .A(\iRF_stage/reg_bank/reg_bank[958] ), .B(n11), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1096 ) );
  MX2X1 U1466 ( .A(\iRF_stage/reg_bank/reg_bank[957] ), .B(n13), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1095 ) );
  MX2X1 U1467 ( .A(\iRF_stage/reg_bank/reg_bank[956] ), .B(n14), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1094 ) );
  MX2X1 U1468 ( .A(\iRF_stage/reg_bank/reg_bank[955] ), .B(n15), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1093 ) );
  MX2X1 U1469 ( .A(\iRF_stage/reg_bank/reg_bank[954] ), .B(n16), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1092 ) );
  MX2X1 U1470 ( .A(\iRF_stage/reg_bank/reg_bank[953] ), .B(n17), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1091 ) );
  MX2X1 U1471 ( .A(\iRF_stage/reg_bank/reg_bank[952] ), .B(n18), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1090 ) );
  MX2X1 U1472 ( .A(\iRF_stage/reg_bank/reg_bank[951] ), .B(n19), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1089 ) );
  MX2X1 U1473 ( .A(\iRF_stage/reg_bank/reg_bank[950] ), .B(n20), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1088 ) );
  MX2X1 U1474 ( .A(\iRF_stage/reg_bank/reg_bank[949] ), .B(n21), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1087 ) );
  MX2X1 U1475 ( .A(\iRF_stage/reg_bank/reg_bank[948] ), .B(n22), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1086 ) );
  MX2X1 U1476 ( .A(\iRF_stage/reg_bank/reg_bank[947] ), .B(n24), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1085 ) );
  MX2X1 U1477 ( .A(\iRF_stage/reg_bank/reg_bank[946] ), .B(n25), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1084 ) );
  MX2X1 U1478 ( .A(\iRF_stage/reg_bank/reg_bank[945] ), .B(n26), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1083 ) );
  MX2X1 U1479 ( .A(\iRF_stage/reg_bank/reg_bank[944] ), .B(n27), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1082 ) );
  MX2X1 U1480 ( .A(\iRF_stage/reg_bank/reg_bank[943] ), .B(n28), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1081 ) );
  MX2X1 U1481 ( .A(\iRF_stage/reg_bank/reg_bank[942] ), .B(n29), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1080 ) );
  MX2X1 U1482 ( .A(\iRF_stage/reg_bank/reg_bank[941] ), .B(n30), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1079 ) );
  MX2X1 U1483 ( .A(\iRF_stage/reg_bank/reg_bank[940] ), .B(n31), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1078 ) );
  MX2X1 U1484 ( .A(\iRF_stage/reg_bank/reg_bank[939] ), .B(n32), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1077 ) );
  MX2X1 U1485 ( .A(\iRF_stage/reg_bank/reg_bank[938] ), .B(n33), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1076 ) );
  MX2X1 U1486 ( .A(\iRF_stage/reg_bank/reg_bank[937] ), .B(n3), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1075 ) );
  MX2X1 U1487 ( .A(\iRF_stage/reg_bank/reg_bank[936] ), .B(n4), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1074 ) );
  MX2X1 U1488 ( .A(\iRF_stage/reg_bank/reg_bank[935] ), .B(n5), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1073 ) );
  MX2X1 U1489 ( .A(\iRF_stage/reg_bank/reg_bank[934] ), .B(n6), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1072 ) );
  MX2X1 U1490 ( .A(\iRF_stage/reg_bank/reg_bank[933] ), .B(n7), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1071 ) );
  MX2X1 U1491 ( .A(\iRF_stage/reg_bank/reg_bank[932] ), .B(n8), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1070 ) );
  MX2X1 U1492 ( .A(\iRF_stage/reg_bank/reg_bank[931] ), .B(n9), .S0(n645), .Y(
        \iRF_stage/reg_bank/n1069 ) );
  MX2X1 U1493 ( .A(\iRF_stage/reg_bank/reg_bank[930] ), .B(n12), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1068 ) );
  MX2X1 U1494 ( .A(\iRF_stage/reg_bank/reg_bank[929] ), .B(n23), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1067 ) );
  MX2X1 U1495 ( .A(\iRF_stage/reg_bank/reg_bank[928] ), .B(n34), .S0(n645), 
        .Y(\iRF_stage/reg_bank/n1066 ) );
  AND2X1 U1496 ( .A(n611), .B(n602), .Y(n645) );
  NOR3X1 U1497 ( .A(\iRF_stage/reg_bank/r_wraddress[0] ), .B(
        \iRF_stage/reg_bank/r_wraddress[2] ), .C(n639), .Y(n611) );
  MX2X1 U1498 ( .A(\iRF_stage/reg_bank/reg_bank[927] ), .B(n10), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1065 ) );
  MX2X1 U1499 ( .A(\iRF_stage/reg_bank/reg_bank[926] ), .B(n11), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1064 ) );
  MX2X1 U1500 ( .A(\iRF_stage/reg_bank/reg_bank[925] ), .B(n13), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1063 ) );
  MX2X1 U1501 ( .A(\iRF_stage/reg_bank/reg_bank[924] ), .B(n14), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1062 ) );
  MX2X1 U1502 ( .A(\iRF_stage/reg_bank/reg_bank[923] ), .B(n15), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1061 ) );
  MX2X1 U1503 ( .A(\iRF_stage/reg_bank/reg_bank[922] ), .B(n16), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1060 ) );
  MX2X1 U1504 ( .A(\iRF_stage/reg_bank/reg_bank[921] ), .B(n17), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1059 ) );
  MX2X1 U1505 ( .A(\iRF_stage/reg_bank/reg_bank[920] ), .B(n18), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1058 ) );
  MX2X1 U1506 ( .A(\iRF_stage/reg_bank/reg_bank[919] ), .B(n19), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1057 ) );
  MX2X1 U1507 ( .A(\iRF_stage/reg_bank/reg_bank[918] ), .B(n20), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1056 ) );
  MX2X1 U1508 ( .A(\iRF_stage/reg_bank/reg_bank[917] ), .B(n21), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1055 ) );
  MX2X1 U1509 ( .A(\iRF_stage/reg_bank/reg_bank[916] ), .B(n22), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1054 ) );
  MX2X1 U1510 ( .A(\iRF_stage/reg_bank/reg_bank[915] ), .B(n24), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1053 ) );
  MX2X1 U1511 ( .A(\iRF_stage/reg_bank/reg_bank[914] ), .B(n25), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1052 ) );
  MX2X1 U1512 ( .A(\iRF_stage/reg_bank/reg_bank[913] ), .B(n26), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1051 ) );
  MX2X1 U1513 ( .A(\iRF_stage/reg_bank/reg_bank[912] ), .B(n27), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1050 ) );
  MX2X1 U1514 ( .A(\iRF_stage/reg_bank/reg_bank[911] ), .B(n28), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1049 ) );
  MX2X1 U1515 ( .A(\iRF_stage/reg_bank/reg_bank[910] ), .B(n29), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1048 ) );
  MX2X1 U1516 ( .A(\iRF_stage/reg_bank/reg_bank[909] ), .B(n30), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1047 ) );
  MX2X1 U1517 ( .A(\iRF_stage/reg_bank/reg_bank[908] ), .B(n31), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1046 ) );
  MX2X1 U1518 ( .A(\iRF_stage/reg_bank/reg_bank[907] ), .B(n32), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1045 ) );
  MX2X1 U1519 ( .A(\iRF_stage/reg_bank/reg_bank[906] ), .B(n33), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1044 ) );
  MX2X1 U1520 ( .A(\iRF_stage/reg_bank/reg_bank[905] ), .B(n3), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1043 ) );
  MX2X1 U1521 ( .A(\iRF_stage/reg_bank/reg_bank[904] ), .B(n4), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1042 ) );
  MX2X1 U1522 ( .A(\iRF_stage/reg_bank/reg_bank[903] ), .B(n5), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1041 ) );
  MX2X1 U1523 ( .A(\iRF_stage/reg_bank/reg_bank[902] ), .B(n6), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1040 ) );
  MX2X1 U1524 ( .A(\iRF_stage/reg_bank/reg_bank[901] ), .B(n7), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1039 ) );
  MX2X1 U1525 ( .A(\iRF_stage/reg_bank/reg_bank[900] ), .B(n8), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1038 ) );
  MX2X1 U1526 ( .A(\iRF_stage/reg_bank/reg_bank[899] ), .B(n9), .S0(n646), .Y(
        \iRF_stage/reg_bank/n1037 ) );
  MX2X1 U1527 ( .A(\iRF_stage/reg_bank/reg_bank[898] ), .B(n12), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1036 ) );
  MX2X1 U1528 ( .A(\iRF_stage/reg_bank/reg_bank[897] ), .B(n23), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1035 ) );
  MX2X1 U1529 ( .A(\iRF_stage/reg_bank/reg_bank[896] ), .B(n34), .S0(n646), 
        .Y(\iRF_stage/reg_bank/n1034 ) );
  AND2X1 U1530 ( .A(n613), .B(n602), .Y(n646) );
  NOR3X1 U1531 ( .A(n639), .B(\iRF_stage/reg_bank/r_wraddress[2] ), .C(n642), 
        .Y(n613) );
  MX2X1 U1532 ( .A(\iRF_stage/reg_bank/reg_bank[895] ), .B(n10), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1033 ) );
  MX2X1 U1533 ( .A(\iRF_stage/reg_bank/reg_bank[894] ), .B(n11), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1032 ) );
  MX2X1 U1534 ( .A(\iRF_stage/reg_bank/reg_bank[893] ), .B(n13), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1031 ) );
  MX2X1 U1535 ( .A(\iRF_stage/reg_bank/reg_bank[892] ), .B(n14), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1030 ) );
  MX2X1 U1536 ( .A(\iRF_stage/reg_bank/reg_bank[891] ), .B(n15), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1029 ) );
  MX2X1 U1537 ( .A(\iRF_stage/reg_bank/reg_bank[890] ), .B(n16), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1028 ) );
  MX2X1 U1538 ( .A(\iRF_stage/reg_bank/reg_bank[889] ), .B(n17), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1027 ) );
  MX2X1 U1539 ( .A(\iRF_stage/reg_bank/reg_bank[888] ), .B(n18), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1026 ) );
  MX2X1 U1540 ( .A(\iRF_stage/reg_bank/reg_bank[887] ), .B(n19), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1025 ) );
  MX2X1 U1541 ( .A(\iRF_stage/reg_bank/reg_bank[886] ), .B(n20), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1024 ) );
  MX2X1 U1542 ( .A(\iRF_stage/reg_bank/reg_bank[885] ), .B(n21), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1023 ) );
  MX2X1 U1543 ( .A(\iRF_stage/reg_bank/reg_bank[884] ), .B(n22), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1022 ) );
  MX2X1 U1544 ( .A(\iRF_stage/reg_bank/reg_bank[883] ), .B(n24), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1021 ) );
  MX2X1 U1545 ( .A(\iRF_stage/reg_bank/reg_bank[882] ), .B(n25), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1020 ) );
  MX2X1 U1546 ( .A(\iRF_stage/reg_bank/reg_bank[881] ), .B(n26), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1019 ) );
  MX2X1 U1547 ( .A(\iRF_stage/reg_bank/reg_bank[880] ), .B(n27), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1018 ) );
  MX2X1 U1548 ( .A(\iRF_stage/reg_bank/reg_bank[879] ), .B(n28), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1017 ) );
  MX2X1 U1549 ( .A(\iRF_stage/reg_bank/reg_bank[878] ), .B(n29), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1016 ) );
  MX2X1 U1550 ( .A(\iRF_stage/reg_bank/reg_bank[877] ), .B(n30), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1015 ) );
  MX2X1 U1551 ( .A(\iRF_stage/reg_bank/reg_bank[876] ), .B(n31), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1014 ) );
  MX2X1 U1552 ( .A(\iRF_stage/reg_bank/reg_bank[875] ), .B(n32), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1013 ) );
  MX2X1 U1553 ( .A(\iRF_stage/reg_bank/reg_bank[874] ), .B(n33), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1012 ) );
  MX2X1 U1554 ( .A(\iRF_stage/reg_bank/reg_bank[873] ), .B(n3), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1011 ) );
  MX2X1 U1555 ( .A(\iRF_stage/reg_bank/reg_bank[872] ), .B(n4), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1010 ) );
  MX2X1 U1556 ( .A(\iRF_stage/reg_bank/reg_bank[871] ), .B(n5), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1009 ) );
  MX2X1 U1557 ( .A(\iRF_stage/reg_bank/reg_bank[870] ), .B(n6), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1008 ) );
  MX2X1 U1558 ( .A(\iRF_stage/reg_bank/reg_bank[869] ), .B(n7), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1007 ) );
  MX2X1 U1559 ( .A(\iRF_stage/reg_bank/reg_bank[868] ), .B(n8), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1006 ) );
  MX2X1 U1560 ( .A(\iRF_stage/reg_bank/reg_bank[867] ), .B(n9), .S0(n647), .Y(
        \iRF_stage/reg_bank/n1005 ) );
  MX2X1 U1561 ( .A(\iRF_stage/reg_bank/reg_bank[866] ), .B(n12), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1004 ) );
  MX2X1 U1562 ( .A(\iRF_stage/reg_bank/reg_bank[865] ), .B(n23), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1003 ) );
  MX2X1 U1563 ( .A(\iRF_stage/reg_bank/reg_bank[864] ), .B(n34), .S0(n647), 
        .Y(\iRF_stage/reg_bank/n1002 ) );
  AND2X1 U1564 ( .A(n615), .B(n602), .Y(n647) );
  NOR3X1 U1565 ( .A(\iRF_stage/reg_bank/r_wraddress[0] ), .B(
        \iRF_stage/reg_bank/r_wraddress[1] ), .C(n640), .Y(n615) );
  MX2X1 U1566 ( .A(\iRF_stage/reg_bank/reg_bank[863] ), .B(n10), .S0(n599), 
        .Y(\iRF_stage/reg_bank/n1001 ) );
  MX2X1 U1567 ( .A(\iRF_stage/reg_bank/reg_bank[862] ), .B(n11), .S0(n599), 
        .Y(\iRF_stage/reg_bank/n1000 ) );
  AND2X1 U1568 ( .A(n617), .B(n602), .Y(n599) );
  NOR3BX1 U1569 ( .AN(\iRF_stage/reg_bank/r_wren ), .B(
        \iRF_stage/reg_bank/r_wraddress[3] ), .C(
        \iRF_stage/reg_bank/r_wraddress[4] ), .Y(n602) );
  NOR3X1 U1570 ( .A(n642), .B(\iRF_stage/reg_bank/r_wraddress[1] ), .C(n640), 
        .Y(n617) );
  CLKINVX1 U1571 ( .A(\iRF_stage/reg_bank/r_wraddress[2] ), .Y(n640) );
  NOR3X1 U1572 ( .A(n648), .B(\iRF_stage/MAIN_FSM/CurrState[0] ), .C(n649), 
        .Y(\iRF_stage/MAIN_FSM/n57 ) );
  OAI2BB1X1 U1573 ( .A0N(n466), .A1N(n650), .B0(rst), .Y(
        \iRF_stage/MAIN_FSM/N52 ) );
  OAI211X1 U1574 ( .A0(n649), .A1(n651), .B0(n652), .C0(rst), .Y(
        \iRF_stage/MAIN_FSM/N51 ) );
  CLKINVX1 U1575 ( .A(n653), .Y(n652) );
  AOI31X1 U1576 ( .A0(n654), .A1(n655), .A2(n656), .B0(n535), .Y(n653) );
  CLKINVX1 U1577 ( .A(n466), .Y(n535) );
  NAND2X1 U1578 ( .A(n657), .B(n658), .Y(n466) );
  NAND2X1 U1579 ( .A(n659), .B(n660), .Y(n651) );
  AOI31X1 U1580 ( .A0(n661), .A1(n662), .A2(n663), .B0(n648), .Y(
        \iRF_stage/MAIN_FSM/N50 ) );
  CLKINVX1 U1581 ( .A(rst), .Y(n648) );
  AOI31X1 U1582 ( .A0(\iRF_stage/MAIN_FSM/CurrState[1] ), .A1(n660), .A2(n664), 
        .B0(n665), .Y(n663) );
  XOR2X1 U1583 ( .A(n37), .B(n666), .Y(n665) );
  NOR2X1 U1584 ( .A(\iRF_stage/MAIN_FSM/CurrState[0] ), .B(
        \iRF_stage/MAIN_FSM/CurrState[1] ), .Y(n666) );
  CLKINVX1 U1585 ( .A(n659), .Y(n664) );
  NAND4X1 U1586 ( .A(n1937), .B(n41), .C(n306), .D(n667), .Y(n659) );
  NOR3X1 U1587 ( .A(\iRF_stage/MAIN_FSM/delay_counter[1] ), .B(
        \iRF_stage/MAIN_FSM/delay_counter[3] ), .C(
        \iRF_stage/MAIN_FSM/delay_counter[2] ), .Y(n667) );
  OR3X1 U1588 ( .A(n658), .B(n668), .C(n669), .Y(n662) );
  NAND2X1 U1589 ( .A(n670), .B(n37), .Y(n658) );
  AOI31X1 U1590 ( .A0(n655), .A1(n536), .A2(n671), .B0(
        \iRF_stage/MAIN_FSM/CurrState[2] ), .Y(n661) );
  NOR2X1 U1591 ( .A(n650), .B(n657), .Y(n671) );
  OR4X1 U1592 ( .A(\iRF_stage/MAIN_FSM/CurrState[1] ), .B(n37), .C(n660), .D(
        \iRF_stage/MAIN_FSM/CurrState[2] ), .Y(n657) );
  NOR2X1 U1593 ( .A(n669), .B(n672), .Y(n650) );
  NAND2X1 U1594 ( .A(n669), .B(n668), .Y(n536) );
  NAND2X1 U1595 ( .A(n672), .B(n669), .Y(n655) );
  NAND3X1 U1596 ( .A(n673), .B(n674), .C(n675), .Y(n669) );
  CLKINVX1 U1597 ( .A(n668), .Y(n672) );
  OAI211X1 U1598 ( .A0(n676), .A1(n677), .B0(n673), .C0(n674), .Y(n668) );
  XOR2X1 U1599 ( .A(n41), .B(\iRF_stage/MAIN_FSM/add_58/carry[5] ), .Y(
        \iRF_stage/MAIN_FSM/N37 ) );
  MXI2X1 U1600 ( .A(n678), .B(n679), .S0(n284), .Y(dout[9]) );
  MXI2X1 U1601 ( .A(n680), .B(n681), .S0(n284), .Y(dout[8]) );
  OAI222X1 U1602 ( .A0(n283), .A1(n682), .B0(n683), .B1(n684), .C0(n685), .C1(
        BUS5985[2]), .Y(dout[31]) );
  CLKINVX1 U1603 ( .A(BUS9884[31]), .Y(n683) );
  OAI222X1 U1604 ( .A0(n283), .A1(n686), .B0(n687), .B1(n684), .C0(n688), .C1(
        BUS5985[2]), .Y(dout[30]) );
  CLKINVX1 U1605 ( .A(BUS9884[30]), .Y(n687) );
  OAI222X1 U1606 ( .A0(n283), .A1(n689), .B0(n690), .B1(n684), .C0(n691), .C1(
        BUS5985[2]), .Y(dout[29]) );
  CLKINVX1 U1607 ( .A(BUS9884[29]), .Y(n690) );
  OAI222X1 U1608 ( .A0(n283), .A1(n692), .B0(n693), .B1(n684), .C0(n694), .C1(
        BUS5985[2]), .Y(dout[28]) );
  CLKINVX1 U1609 ( .A(BUS9884[28]), .Y(n693) );
  OAI222X1 U1610 ( .A0(n283), .A1(n695), .B0(n696), .B1(n684), .C0(n697), .C1(
        BUS5985[2]), .Y(dout[27]) );
  CLKINVX1 U1611 ( .A(BUS9884[27]), .Y(n696) );
  OAI222X1 U1612 ( .A0(n283), .A1(n698), .B0(n699), .B1(n684), .C0(n700), .C1(
        BUS5985[2]), .Y(dout[26]) );
  CLKINVX1 U1613 ( .A(BUS9884[26]), .Y(n699) );
  OAI222X1 U1614 ( .A0(n283), .A1(n678), .B0(n701), .B1(n684), .C0(n679), .C1(
        BUS5985[2]), .Y(dout[25]) );
  CLKINVX1 U1615 ( .A(BUS9884[25]), .Y(n701) );
  CLKINVX1 U1616 ( .A(BUS9884[9]), .Y(n678) );
  OAI222X1 U1617 ( .A0(n283), .A1(n680), .B0(n702), .B1(n684), .C0(n681), .C1(
        BUS5985[2]), .Y(dout[24]) );
  CLKINVX1 U1618 ( .A(BUS9884[24]), .Y(n702) );
  CLKINVX1 U1619 ( .A(BUS9884[8]), .Y(n680) );
  OAI22X1 U1620 ( .A0(n685), .A1(n703), .B0(n704), .B1(n684), .Y(dout[23]) );
  CLKINVX1 U1621 ( .A(BUS9884[23]), .Y(n704) );
  OAI22X1 U1622 ( .A0(n688), .A1(n703), .B0(n705), .B1(n684), .Y(dout[22]) );
  CLKINVX1 U1623 ( .A(BUS9884[22]), .Y(n705) );
  OAI22X1 U1624 ( .A0(n691), .A1(n703), .B0(n706), .B1(n684), .Y(dout[21]) );
  CLKINVX1 U1625 ( .A(BUS9884[21]), .Y(n706) );
  OAI22X1 U1626 ( .A0(n694), .A1(n703), .B0(n707), .B1(n684), .Y(dout[20]) );
  CLKINVX1 U1627 ( .A(BUS9884[20]), .Y(n707) );
  OAI22X1 U1628 ( .A0(n697), .A1(n703), .B0(n708), .B1(n684), .Y(dout[19]) );
  CLKINVX1 U1629 ( .A(BUS9884[19]), .Y(n708) );
  OAI22X1 U1630 ( .A0(n700), .A1(n703), .B0(n709), .B1(n684), .Y(dout[18]) );
  CLKINVX1 U1631 ( .A(BUS9884[18]), .Y(n709) );
  OAI22X1 U1632 ( .A0(n679), .A1(n703), .B0(n710), .B1(n684), .Y(dout[17]) );
  CLKINVX1 U1633 ( .A(BUS9884[17]), .Y(n710) );
  CLKINVX1 U1634 ( .A(dout[1]), .Y(n679) );
  OAI222X1 U1635 ( .A0(n711), .A1(n712), .B0(n713), .B1(n714), .C0(n715), .C1(
        n716), .Y(dout[1]) );
  OAI22X1 U1636 ( .A0(n681), .A1(n703), .B0(n717), .B1(n684), .Y(dout[16]) );
  CLKINVX1 U1637 ( .A(BUS9884[16]), .Y(n717) );
  OAI21X1 U1638 ( .A0(BUS5985[2]), .A1(n283), .B0(n684), .Y(n703) );
  NAND2X1 U1639 ( .A(n283), .B(BUS5985[2]), .Y(n684) );
  CLKINVX1 U1640 ( .A(dout[0]), .Y(n681) );
  MXI2X1 U1641 ( .A(n682), .B(n685), .S0(n284), .Y(dout[15]) );
  CLKINVX1 U1642 ( .A(dout[7]), .Y(n685) );
  OAI222X1 U1643 ( .A0(n711), .A1(n718), .B0(n719), .B1(n714), .C0(n715), .C1(
        n720), .Y(dout[7]) );
  CLKINVX1 U1644 ( .A(BUS9884[15]), .Y(n682) );
  MXI2X1 U1645 ( .A(n686), .B(n688), .S0(n284), .Y(dout[14]) );
  CLKINVX1 U1646 ( .A(dout[6]), .Y(n688) );
  OAI222X1 U1647 ( .A0(n711), .A1(n721), .B0(n722), .B1(n714), .C0(n715), .C1(
        n723), .Y(dout[6]) );
  CLKINVX1 U1648 ( .A(BUS9884[14]), .Y(n686) );
  MXI2X1 U1649 ( .A(n689), .B(n691), .S0(n284), .Y(dout[13]) );
  CLKINVX1 U1650 ( .A(dout[5]), .Y(n691) );
  OAI222X1 U1651 ( .A0(n711), .A1(n724), .B0(n725), .B1(n714), .C0(n715), .C1(
        n726), .Y(dout[5]) );
  CLKINVX1 U1652 ( .A(BUS9884[13]), .Y(n689) );
  MXI2X1 U1653 ( .A(n692), .B(n694), .S0(n284), .Y(dout[12]) );
  CLKINVX1 U1654 ( .A(dout[4]), .Y(n694) );
  OAI222X1 U1655 ( .A0(n711), .A1(n727), .B0(n728), .B1(n714), .C0(n715), .C1(
        n729), .Y(dout[4]) );
  CLKINVX1 U1656 ( .A(BUS9884[12]), .Y(n692) );
  MXI2X1 U1657 ( .A(n695), .B(n697), .S0(n284), .Y(dout[11]) );
  CLKINVX1 U1658 ( .A(dout[3]), .Y(n697) );
  OAI222X1 U1659 ( .A0(n711), .A1(n730), .B0(n731), .B1(n714), .C0(n715), .C1(
        n732), .Y(dout[3]) );
  CLKINVX1 U1660 ( .A(BUS9884[11]), .Y(n695) );
  MXI2X1 U1661 ( .A(n698), .B(n700), .S0(n284), .Y(dout[10]) );
  CLKINVX1 U1662 ( .A(dout[2]), .Y(n700) );
  OAI222X1 U1663 ( .A0(n711), .A1(n733), .B0(n734), .B1(n714), .C0(n715), .C1(
        n735), .Y(dout[2]) );
  CLKINVX1 U1664 ( .A(BUS9884[10]), .Y(n698) );
  OAI222X1 U1665 ( .A0(n711), .A1(n736), .B0(n737), .B1(n714), .C0(n715), .C1(
        n738), .Y(dout[0]) );
  OAI2BB2X1 U1666 ( .B0(n739), .B1(n740), .A0N(
        \decoder_pipe/pipereg/BUS4987[0] ), .A1N(n538), .Y(
        \decoder_pipe/pipereg/U6/n4 ) );
  AOI211X1 U1667 ( .A0(n741), .A1(n742), .B0(n743), .C0(
        \decoder_pipe/BUS2110[0] ), .Y(n739) );
  OAI2BB2X1 U1668 ( .B0(n744), .B1(n740), .A0N(
        \decoder_pipe/pipereg/BUS5639[0] ), .A1N(n538), .Y(
        \decoder_pipe/pipereg/U11/n4 ) );
  OAI2BB2X1 U1669 ( .B0(n745), .B1(n740), .A0N(
        \decoder_pipe/pipereg/BUS5651[0] ), .A1N(n538), .Y(
        \decoder_pipe/pipereg/U10/n4 ) );
  NOR2X1 U1670 ( .A(n649), .B(n660), .Y(n538) );
  OR2X1 U1671 ( .A(n459), .B(\iRF_stage/MAIN_FSM/CurrState[2] ), .Y(n649) );
  NOR2BX1 U1672 ( .AN(n746), .B(n467), .Y(n1933) );
  OAI211X1 U1673 ( .A0(n458), .A1(n459), .B0(n598), .C0(n747), .Y(n467) );
  XOR2X1 U1674 ( .A(\iRF_stage/MAIN_FSM/n17 ), .B(n670), .Y(n747) );
  NOR3X1 U1675 ( .A(\iRF_stage/MAIN_FSM/CurrState[1] ), .B(
        \iRF_stage/MAIN_FSM/CurrState[2] ), .C(
        \iRF_stage/MAIN_FSM/CurrState[0] ), .Y(n670) );
  NAND2X1 U1676 ( .A(n1935), .B(\iRF_stage/MAIN_FSM/CurrState[0] ), .Y(n598)
         );
  NOR3X1 U1677 ( .A(n37), .B(\iRF_stage/MAIN_FSM/CurrState[1] ), .C(n748), .Y(
        n1935) );
  NAND2X1 U1678 ( .A(\iRF_stage/MAIN_FSM/CurrState[1] ), .B(
        \iRF_stage/MAIN_FSM/n17 ), .Y(n459) );
  NAND2X1 U1679 ( .A(\iRF_stage/MAIN_FSM/CurrState[2] ), .B(n660), .Y(n458) );
  CLKINVX1 U1680 ( .A(\iRF_stage/MAIN_FSM/CurrState[0] ), .Y(n660) );
  OAI2BB1X1 U1681 ( .A0N(\iRF_stage/MAIN_FSM/CurrState[0] ), .A1N(n748), .B0(
        \iRF_stage/MAIN_FSM/CurrState[1] ), .Y(n746) );
  CLKINVX1 U1682 ( .A(\iRF_stage/MAIN_FSM/CurrState[2] ), .Y(n748) );
  OR2X1 U1683 ( .A(NET767), .B(\decoder_pipe/pipereg/BUS7822[0] ), .Y(
        \decoder_pipe/pipereg/NET7643 ) );
  OAI211X1 U1684 ( .A0(n749), .A1(n750), .B0(n674), .C0(n751), .Y(
        \decoder_pipe/BUS2110[1] ) );
  NAND4X1 U1685 ( .A(n674), .B(n752), .C(n753), .D(n754), .Y(
        \decoder_pipe/BUS2110[0] ) );
  AOI2BB2X1 U1686 ( .B0(n755), .B1(n756), .A0N(n757), .A1N(n758), .Y(n754) );
  NAND3X1 U1687 ( .A(n751), .B(n654), .C(n759), .Y(\decoder_pipe/BUS2102[2] )
         );
  AOI211X1 U1688 ( .A0(n760), .A1(n761), .B0(n762), .C0(n763), .Y(n759) );
  OAI21X1 U1689 ( .A0(n676), .A1(n677), .B0(n656), .Y(
        \decoder_pipe/BUS2102[1] ) );
  NAND4X1 U1690 ( .A(n764), .B(n765), .C(n760), .D(n766), .Y(n656) );
  NOR2X1 U1691 ( .A(n767), .B(n758), .Y(n766) );
  NAND4X1 U1692 ( .A(n537), .B(n768), .C(n769), .D(n770), .Y(
        \decoder_pipe/BUS2102[0] ) );
  AOI21X1 U1693 ( .A0(n760), .A1(n761), .B0(n771), .Y(n770) );
  NAND2X1 U1694 ( .A(n772), .B(n773), .Y(n761) );
  NOR2X1 U1695 ( .A(n774), .B(n775), .Y(n537) );
  NAND2X1 U1696 ( .A(n751), .B(n768), .Y(\decoder_pipe/BUS2094[1] ) );
  OAI211X1 U1697 ( .A0(n776), .A1(n772), .B0(n675), .C0(n674), .Y(
        \decoder_pipe/BUS2094[0] ) );
  OAI211X1 U1698 ( .A0(n776), .A1(n772), .B0(n751), .C0(n777), .Y(
        \decoder_pipe/BUS2086[1] ) );
  NOR2X1 U1699 ( .A(n778), .B(n743), .Y(n751) );
  OAI221X1 U1700 ( .A0(n779), .A1(n780), .B0(n781), .B1(n749), .C0(n782), .Y(
        n743) );
  OAI221X1 U1701 ( .A0(n783), .A1(n756), .B0(n784), .B1(n767), .C0(n765), .Y(
        n772) );
  NOR2X1 U1702 ( .A(n785), .B(n764), .Y(n784) );
  OAI2BB1X1 U1703 ( .A0N(ins_i[1]), .A1N(n786), .B0(n787), .Y(n756) );
  NAND3X1 U1704 ( .A(n788), .B(n782), .C(n654), .Y(\decoder_pipe/BUS2072[2] )
         );
  AOI221XL U1705 ( .A0(n789), .A1(n790), .B0(n791), .B1(n741), .C0(
        \decoder_pipe/BUS2056[2] ), .Y(n654) );
  NAND4BX1 U1706 ( .AN(n792), .B(n793), .C(n794), .D(n795), .Y(
        \decoder_pipe/BUS2072[0] ) );
  NOR2X1 U1707 ( .A(\decoder_pipe/BUS2086[0] ), .B(n775), .Y(n794) );
  CLKINVX1 U1708 ( .A(n673), .Y(n775) );
  NAND2X1 U1709 ( .A(n796), .B(n791), .Y(n673) );
  NAND2X1 U1710 ( .A(n674), .B(n788), .Y(\decoder_pipe/BUS2086[0] ) );
  NAND4X1 U1711 ( .A(n755), .B(n797), .C(n786), .D(n787), .Y(n788) );
  NAND2X1 U1712 ( .A(ins_i[0]), .B(n764), .Y(n797) );
  OAI221X1 U1713 ( .A0(n798), .A1(n799), .B0(n779), .B1(n750), .C0(n800), .Y(
        \decoder_pipe/BUS2064[2] ) );
  CLKINVX1 U1714 ( .A(n801), .Y(n799) );
  NAND4X1 U1715 ( .A(n802), .B(n752), .C(n800), .D(n803), .Y(
        \decoder_pipe/BUS2064[1] ) );
  AOI22X1 U1716 ( .A0(n801), .A1(n798), .B0(n804), .B1(n805), .Y(n803) );
  OAI22X1 U1717 ( .A0(n806), .A1(n807), .B0(n808), .B1(n809), .Y(
        \decoder_pipe/BUS2056[2] ) );
  OAI22X1 U1718 ( .A0(n806), .A1(n810), .B0(n811), .B1(n808), .Y(
        \decoder_pipe/BUS2056[1] ) );
  AOI2BB1X1 U1719 ( .A0N(\iRF_stage/BUS3236[0] ), .A1N(n809), .B0(n812), .Y(
        n811) );
  NAND3BX1 U1720 ( .AN(\iRF_stage/BUS3236[1] ), .B(n813), .C(n814), .Y(n809)
         );
  NOR3X1 U1721 ( .A(\iRF_stage/BUS3236[2] ), .B(\iRF_stage/BUS3236[4] ), .C(
        \iRF_stage/BUS3236[3] ), .Y(n814) );
  OAI22X1 U1722 ( .A0(n808), .A1(n810), .B0(n781), .B1(n806), .Y(
        \decoder_pipe/BUS2056[0] ) );
  CLKINVX1 U1723 ( .A(n791), .Y(n806) );
  CLKINVX1 U1724 ( .A(n789), .Y(n781) );
  NAND4X1 U1725 ( .A(n752), .B(n815), .C(n769), .D(n816), .Y(
        \decoder_pipe/BUS2040[4] ) );
  AOI221XL U1726 ( .A0(n817), .A1(ins_i[3]), .B0(ins_i[2]), .B1(n818), .C0(
        n774), .Y(n816) );
  OAI211X1 U1727 ( .A0(n749), .A1(n807), .B0(n819), .C0(n820), .Y(n774) );
  AOI2BB2X1 U1728 ( .B0(n742), .B1(n813), .A0N(n810), .A1N(n779), .Y(n820) );
  CLKINVX1 U1729 ( .A(n821), .Y(n818) );
  CLKINVX1 U1730 ( .A(n753), .Y(n817) );
  OAI211X1 U1731 ( .A0(ins_i[2]), .A1(n821), .B0(n793), .C0(n777), .Y(
        \decoder_pipe/BUS2040[3] ) );
  NOR3BX1 U1732 ( .AN(n815), .B(n822), .C(n762), .Y(n777) );
  CLKINVX1 U1733 ( .A(n771), .Y(n793) );
  OAI21X1 U1734 ( .A0(n780), .A1(n749), .B0(n745), .Y(n771) );
  NAND4BX1 U1735 ( .AN(n823), .B(n824), .C(n768), .D(n825), .Y(
        \decoder_pipe/BUS2040[2] ) );
  NAND2X1 U1736 ( .A(ins_i[1]), .B(n826), .Y(n825) );
  OAI31X1 U1737 ( .A0(n827), .A1(ins_i[2]), .A2(n828), .B0(n821), .Y(n826) );
  CLKINVX1 U1738 ( .A(n1928), .Y(n768) );
  NAND2X1 U1739 ( .A(n795), .B(n752), .Y(n1928) );
  CLKINVX1 U1740 ( .A(n762), .Y(n795) );
  OAI32X1 U1741 ( .A0(n829), .A1(ins_i[28]), .A2(n749), .B0(n779), .B1(n750), 
        .Y(n762) );
  NOR2X1 U1742 ( .A(n805), .B(n742), .Y(n779) );
  OAI211X1 U1743 ( .A0(n749), .A1(n780), .B0(n744), .C0(n819), .Y(n823) );
  CLKINVX1 U1744 ( .A(n778), .Y(n744) );
  OAI2BB1X1 U1745 ( .A0N(n742), .A1N(n741), .B0(n745), .Y(n778) );
  NOR3BX1 U1746 ( .AN(n800), .B(n1931), .C(n801), .Y(n745) );
  NOR2X1 U1747 ( .A(n829), .B(n808), .Y(n801) );
  NAND2X1 U1748 ( .A(n830), .B(n831), .Y(n829) );
  OAI21X1 U1749 ( .A0(n808), .A1(n750), .B0(n802), .Y(n1931) );
  NAND4X1 U1750 ( .A(ins_i[28]), .B(ins_i[26]), .C(n830), .D(n790), .Y(n802)
         );
  NAND2X1 U1751 ( .A(n791), .B(n804), .Y(n800) );
  CLKINVX1 U1752 ( .A(n750), .Y(n804) );
  NAND3X1 U1753 ( .A(n830), .B(n798), .C(ins_i[26]), .Y(n750) );
  NOR2X1 U1754 ( .A(n832), .B(ins_i[30]), .Y(n830) );
  NOR2X1 U1755 ( .A(n796), .B(n813), .Y(n780) );
  NAND3X1 U1756 ( .A(n833), .B(n819), .C(n834), .Y(\decoder_pipe/BUS2040[1] )
         );
  AOI211X1 U1757 ( .A0(n805), .A1(n789), .B0(n835), .C0(n836), .Y(n834) );
  CLKINVX1 U1758 ( .A(n752), .Y(n835) );
  NAND2X1 U1759 ( .A(n763), .B(n677), .Y(n752) );
  CLKINVX1 U1760 ( .A(\iRF_stage/BUS3237[2] ), .Y(n677) );
  CLKINVX1 U1761 ( .A(n676), .Y(n763) );
  NAND2X1 U1762 ( .A(n837), .B(n838), .Y(n676) );
  NOR4X1 U1763 ( .A(ins_i[26]), .B(n839), .C(\iRF_stage/BUS3237[4] ), .D(
        \iRF_stage/BUS3237[3] ), .Y(n838) );
  NAND2X1 U1764 ( .A(n798), .B(n832), .Y(n839) );
  CLKINVX1 U1765 ( .A(ins_i[31]), .Y(n832) );
  NOR4BX1 U1766 ( .AN(ins_i[30]), .B(\iRF_stage/BUS3237[1] ), .C(
        \iRF_stage/BUS3237[0] ), .D(n808), .Y(n837) );
  CLKINVX1 U1767 ( .A(n790), .Y(n808) );
  NAND2X1 U1768 ( .A(n810), .B(n807), .Y(n789) );
  AND2X1 U1769 ( .A(n782), .B(n674), .Y(n819) );
  NAND2X1 U1770 ( .A(n813), .B(n791), .Y(n674) );
  NOR2X1 U1771 ( .A(n840), .B(ins_i[29]), .Y(n791) );
  AND3X2 U1772 ( .A(n841), .B(ins_i[26]), .C(n798), .Y(n813) );
  CLKINVX1 U1773 ( .A(ins_i[28]), .Y(n798) );
  MXI2X1 U1774 ( .A(n842), .B(n843), .S0(ins_i[1]), .Y(n833) );
  NAND2X1 U1775 ( .A(n675), .B(n824), .Y(n843) );
  OR2X1 U1776 ( .A(n757), .B(n785), .Y(n824) );
  AOI31X1 U1777 ( .A0(ins_i[5]), .A1(n765), .A2(n786), .B0(n844), .Y(n785) );
  NAND4X1 U1778 ( .A(n782), .B(n815), .C(n845), .D(n846), .Y(
        \decoder_pipe/BUS2040[0] ) );
  AOI221XL U1779 ( .A0(ins_i[1]), .A1(n847), .B0(n741), .B1(n805), .C0(n792), 
        .Y(n846) );
  OAI31X1 U1780 ( .A0(n753), .A1(ins_i[0]), .A2(n767), .B0(n769), .Y(n792) );
  NAND2X1 U1781 ( .A(n742), .B(n796), .Y(n769) );
  NAND4X1 U1782 ( .A(n786), .B(n765), .C(n760), .D(n848), .Y(n753) );
  NOR2X1 U1783 ( .A(n764), .B(n787), .Y(n848) );
  CLKINVX1 U1784 ( .A(n749), .Y(n805) );
  NAND2X1 U1785 ( .A(ins_i[29]), .B(n840), .Y(n749) );
  CLKINVX1 U1786 ( .A(ins_i[27]), .Y(n840) );
  CLKINVX1 U1787 ( .A(n810), .Y(n741) );
  NAND3X1 U1788 ( .A(n841), .B(n831), .C(ins_i[28]), .Y(n810) );
  CLKINVX1 U1789 ( .A(ins_i[26]), .Y(n831) );
  CLKINVX1 U1790 ( .A(n849), .Y(n847) );
  AOI2BB1X1 U1791 ( .A0N(n827), .A1N(n821), .B0(n842), .Y(n849) );
  OAI22X1 U1792 ( .A0(n758), .A1(n828), .B0(n773), .B1(n757), .Y(n842) );
  NAND2X1 U1793 ( .A(n783), .B(n787), .Y(n758) );
  NOR2X1 U1794 ( .A(ins_i[2]), .B(ins_i[0]), .Y(n783) );
  OAI21X1 U1795 ( .A0(n836), .A1(n822), .B0(n827), .Y(n845) );
  CLKINVX1 U1796 ( .A(ins_i[0]), .Y(n827) );
  CLKINVX1 U1797 ( .A(n675), .Y(n822) );
  NAND3X1 U1798 ( .A(n844), .B(n760), .C(ins_i[3]), .Y(n675) );
  NOR3X1 U1799 ( .A(n821), .B(ins_i[1]), .C(n786), .Y(n836) );
  NAND2X1 U1800 ( .A(n755), .B(ins_i[5]), .Y(n821) );
  CLKINVX1 U1801 ( .A(n828), .Y(n755) );
  NAND2X1 U1802 ( .A(n850), .B(n765), .Y(n828) );
  CLKINVX1 U1803 ( .A(ins_i[4]), .Y(n765) );
  NAND4X1 U1804 ( .A(ins_i[0]), .B(n850), .C(n844), .D(n764), .Y(n815) );
  CLKINVX1 U1805 ( .A(ins_i[1]), .Y(n764) );
  CLKINVX1 U1806 ( .A(n773), .Y(n844) );
  NAND3X1 U1807 ( .A(n786), .B(n787), .C(ins_i[4]), .Y(n773) );
  CLKINVX1 U1808 ( .A(ins_i[5]), .Y(n787) );
  CLKINVX1 U1809 ( .A(ins_i[2]), .Y(n786) );
  CLKINVX1 U1810 ( .A(n757), .Y(n850) );
  NAND2X1 U1811 ( .A(n760), .B(n767), .Y(n757) );
  CLKINVX1 U1812 ( .A(ins_i[3]), .Y(n767) );
  CLKINVX1 U1813 ( .A(n776), .Y(n760) );
  NAND2X1 U1814 ( .A(n796), .B(n790), .Y(n776) );
  NOR2X1 U1815 ( .A(ins_i[27]), .B(ins_i[29]), .Y(n790) );
  NOR3BX1 U1816 ( .AN(n841), .B(ins_i[26]), .C(ins_i[28]), .Y(n796) );
  NAND2X1 U1817 ( .A(n812), .B(n742), .Y(n782) );
  AND2X1 U1818 ( .A(ins_i[27]), .B(ins_i[29]), .Y(n742) );
  CLKINVX1 U1819 ( .A(n807), .Y(n812) );
  NAND3X1 U1820 ( .A(n841), .B(ins_i[26]), .C(ins_i[28]), .Y(n807) );
  NOR2X1 U1821 ( .A(ins_i[30]), .B(ins_i[31]), .Y(n841) );
  NAND4X1 U1822 ( .A(n851), .B(n852), .C(n853), .D(n854), .Y(addr_o[9]) );
  AOI221XL U1823 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N185 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N121 ), .B1(n855), .C0(n856), .Y(n854)
         );
  OAI2BB1X1 U1824 ( .A0N(n857), .A1N(\iexec_stage/BUS468[9] ), .B0(n858), .Y(
        n856) );
  MXI2X1 U1825 ( .A(n859), .B(n860), .S0(n568), .Y(n858) );
  NOR2X1 U1826 ( .A(\iexec_stage/BUS468[9] ), .B(n861), .Y(n860) );
  OAI2BB1X1 U1827 ( .A0N(n862), .A1N(\iexec_stage/BUS468[9] ), .B0(n863), .Y(
        n859) );
  AOI22X1 U1828 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N218 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N250 ), .B1(n865), .Y(n853) );
  OAI21X1 U1829 ( .A0(n866), .A1(n867), .B0(n868), .Y(n852) );
  OAI2BB1X1 U1830 ( .A0N(n869), .A1N(n870), .B0(n871), .Y(n851) );
  AOI221XL U1831 ( .A0(n872), .A1(n546), .B0(n873), .B1(n543), .C0(n874), .Y(
        n870) );
  OAI222X1 U1832 ( .A0(n1926), .A1(n875), .B0(n1927), .B1(n876), .C0(n1924), 
        .C1(n877), .Y(n874) );
  AOI221XL U1833 ( .A0(n878), .A1(n539), .B0(n879), .B1(
        \iexec_stage/BUS468[9] ), .C0(n880), .Y(n869) );
  OAI222X1 U1834 ( .A0(n1921), .A1(n881), .B0(n1920), .B1(n882), .C0(n1919), 
        .C1(n883), .Y(n880) );
  NAND4X1 U1835 ( .A(n884), .B(n885), .C(n886), .D(n887), .Y(addr_o[8]) );
  AOI221XL U1836 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N184 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N120 ), .B1(n855), .C0(n888), .Y(n887)
         );
  OAI2BB1X1 U1837 ( .A0N(n539), .A1N(n889), .B0(n890), .Y(n888) );
  MXI2X1 U1838 ( .A(n891), .B(n892), .S0(n569), .Y(n890) );
  NOR2X1 U1839 ( .A(n861), .B(n539), .Y(n892) );
  OAI2BB1X1 U1840 ( .A0N(n862), .A1N(n539), .B0(n863), .Y(n891) );
  AOI22X1 U1841 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N217 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N249 ), .B1(n865), .Y(n886) );
  OAI2BB1X1 U1842 ( .A0N(n893), .A1N(n894), .B0(n868), .Y(n885) );
  OAI2BB1X1 U1843 ( .A0N(n895), .A1N(n896), .B0(n871), .Y(n884) );
  AOI221XL U1844 ( .A0(n897), .A1(n565), .B0(n898), .B1(n546), .C0(n899), .Y(
        n896) );
  OAI22X1 U1845 ( .A0(n1924), .A1(n900), .B0(n1926), .B1(n901), .Y(n899) );
  AOI221XL U1846 ( .A0(n902), .A1(n542), .B0(n903), .B1(n543), .C0(n904), .Y(
        n895) );
  OAI22X1 U1847 ( .A0(n1919), .A1(n905), .B0(n1920), .B1(n883), .Y(n904) );
  NAND4X1 U1848 ( .A(n906), .B(n907), .C(n908), .D(n909), .Y(addr_o[7]) );
  AOI221XL U1849 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N183 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N119 ), .B1(n855), .C0(n910), .Y(n909)
         );
  OAI2BB1X1 U1850 ( .A0N(n540), .A1N(n889), .B0(n911), .Y(n910) );
  MXI2X1 U1851 ( .A(n912), .B(n913), .S0(n570), .Y(n911) );
  NOR2X1 U1852 ( .A(n861), .B(n540), .Y(n913) );
  OAI2BB1X1 U1853 ( .A0N(n862), .A1N(n540), .B0(n863), .Y(n912) );
  AOI22X1 U1854 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N216 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N248 ), .B1(n865), .Y(n908) );
  OAI2BB1X1 U1855 ( .A0N(n914), .A1N(n915), .B0(n868), .Y(n907) );
  OAI2BB1X1 U1856 ( .A0N(n916), .A1N(n917), .B0(n871), .Y(n906) );
  AOI221XL U1857 ( .A0(n898), .A1(\iexec_stage/BUS468[1] ), .B0(n872), .B1(
        n565), .C0(n918), .Y(n917) );
  OAI22X1 U1858 ( .A0(n1922), .A1(n882), .B0(n1925), .B1(n900), .Y(n918) );
  AOI222XL U1859 ( .A0(n878), .A1(n541), .B0(n903), .B1(n544), .C0(n919), .C1(
        n542), .Y(n916) );
  NAND4X1 U1860 ( .A(n920), .B(n921), .C(n922), .D(n923), .Y(addr_o[6]) );
  AOI221XL U1861 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N182 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N118 ), .B1(n855), .C0(n924), .Y(n923)
         );
  OAI2BB1X1 U1862 ( .A0N(n857), .A1N(n541), .B0(n925), .Y(n924) );
  MXI2X1 U1863 ( .A(n926), .B(n927), .S0(n571), .Y(n925) );
  NOR2X1 U1864 ( .A(n861), .B(n541), .Y(n927) );
  OAI2BB1X1 U1865 ( .A0N(n862), .A1N(n541), .B0(n863), .Y(n926) );
  AOI22X1 U1866 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N215 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N247 ), .B1(n865), .Y(n922) );
  OAI2BB1X1 U1867 ( .A0N(n928), .A1N(n929), .B0(n868), .Y(n921) );
  OAI2BB1X1 U1868 ( .A0N(n930), .A1N(n931), .B0(n871), .Y(n920) );
  AOI221XL U1869 ( .A0(n898), .A1(n565), .B0(n873), .B1(
        \iexec_stage/BUS468[1] ), .C0(n932), .Y(n931) );
  OAI22X1 U1870 ( .A0(n1925), .A1(n881), .B0(n1924), .B1(n882), .Y(n932) );
  AOI222XL U1871 ( .A0(n879), .A1(n541), .B0(n919), .B1(n543), .C0(n878), .C1(
        n542), .Y(n930) );
  NAND4X1 U1872 ( .A(n933), .B(n934), .C(n935), .D(n936), .Y(addr_o[5]) );
  AOI221XL U1873 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N181 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N117 ), .B1(n855), .C0(n937), .Y(n936)
         );
  OAI2BB1X1 U1874 ( .A0N(n857), .A1N(n542), .B0(n938), .Y(n937) );
  MXI2X1 U1875 ( .A(n939), .B(n940), .S0(n572), .Y(n938) );
  NOR2X1 U1876 ( .A(n861), .B(n542), .Y(n940) );
  OAI2BB1X1 U1877 ( .A0N(n862), .A1N(n542), .B0(n863), .Y(n939) );
  AOI22X1 U1878 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N214 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N246 ), .B1(n865), .Y(n935) );
  OAI21X1 U1879 ( .A0(n941), .A1(n942), .B0(n868), .Y(n934) );
  OAI2BB1X1 U1880 ( .A0N(n943), .A1N(n944), .B0(n871), .Y(n933) );
  AOI222XL U1881 ( .A0(n903), .A1(\iexec_stage/BUS468[1] ), .B0(n873), .B1(
        n565), .C0(n902), .C1(n546), .Y(n944) );
  AOI222XL U1882 ( .A0(n879), .A1(n542), .B0(n919), .B1(n544), .C0(n878), .C1(
        n543), .Y(n943) );
  NAND4X1 U1883 ( .A(n945), .B(n946), .C(n947), .D(n948), .Y(addr_o[4]) );
  AOI221XL U1884 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N213 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N245 ), .B1(n865), .C0(n949), 
        .Y(n948) );
  OAI22X1 U1885 ( .A0(n950), .A1(n951), .B0(n952), .B1(n953), .Y(n949) );
  NOR2X1 U1886 ( .A(n954), .B(n955), .Y(n952) );
  AOI221XL U1887 ( .A0(n902), .A1(\iexec_stage/BUS468[1] ), .B0(n903), .B1(
        n565), .C0(n956), .Y(n950) );
  OAI22X1 U1888 ( .A0(n1924), .A1(n905), .B0(n1925), .B1(n883), .Y(n956) );
  NAND2X1 U1889 ( .A(n543), .B(n889), .Y(n946) );
  MXI2X1 U1890 ( .A(n957), .B(n958), .S0(n1923), .Y(n945) );
  NOR2X1 U1891 ( .A(n861), .B(n543), .Y(n958) );
  OAI2BB1X1 U1892 ( .A0N(n862), .A1N(n543), .B0(n863), .Y(n957) );
  NAND2X1 U1893 ( .A(n959), .B(n960), .Y(addr_o[3]) );
  AOI221XL U1894 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N212 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N244 ), .B1(n865), .C0(n961), 
        .Y(n960) );
  OAI22X1 U1895 ( .A0(n962), .A1(n951), .B0(n963), .B1(n953), .Y(n961) );
  NOR2X1 U1896 ( .A(n964), .B(n965), .Y(n963) );
  AOI222XL U1897 ( .A0(n878), .A1(n546), .B0(n902), .B1(n565), .C0(n919), .C1(
        \iexec_stage/BUS468[1] ), .Y(n962) );
  AOI221XL U1898 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N179 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N115 ), .B1(n855), .C0(n966), .Y(n959)
         );
  OAI21X1 U1899 ( .A0(n967), .A1(n1924), .B0(n968), .Y(n966) );
  MXI2X1 U1900 ( .A(n969), .B(n970), .S0(n574), .Y(n968) );
  NOR2X1 U1901 ( .A(n861), .B(n544), .Y(n970) );
  OAI2BB1X1 U1902 ( .A0N(n862), .A1N(n544), .B0(n863), .Y(n969) );
  NAND2X1 U1903 ( .A(n971), .B(n972), .Y(addr_o[31]) );
  AOI221XL U1904 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N207 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N208 ), .B1(n871), .C0(n973), .Y(
        n972) );
  AOI221XL U1905 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N143 ), .A1(n855), .B0(
        n974), .B1(\iexec_stage/BUS468[31] ), .C0(n975), .Y(n971) );
  MXI2X1 U1906 ( .A(n976), .B(n977), .S0(n573), .Y(n975) );
  NAND2X1 U1907 ( .A(n978), .B(n1881), .Y(n977) );
  AOI2BB1X1 U1908 ( .A0N(\iexec_stage/BUS468[31] ), .A1N(n953), .B0(n979), .Y(
        n976) );
  OAI211X1 U1909 ( .A0(n980), .A1(n981), .B0(n982), .C0(n983), .Y(n974) );
  MXI2X1 U1910 ( .A(n862), .B(n868), .S0(n573), .Y(n983) );
  CLKINVX1 U1911 ( .A(\iexec_stage/BUS476[31] ), .Y(n573) );
  NAND2X1 U1912 ( .A(n984), .B(n985), .Y(addr_o[30]) );
  AOI221XL U1913 ( .A0(n973), .A1(n986), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N207 ), .B1(n871), .C0(n987), .Y(
        n985) );
  OAI22X1 U1914 ( .A0(n1883), .A1(n988), .B0(n989), .B1(n905), .Y(n987) );
  NOR2X1 U1915 ( .A(n990), .B(n973), .Y(n989) );
  AOI221XL U1916 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N206 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N142 ), .B1(n855), .C0(n991), .Y(n984)
         );
  MXI2X1 U1917 ( .A(n992), .B(n993), .S0(\iexec_stage/BUS476[30] ), .Y(n991)
         );
  NOR2X1 U1918 ( .A(n979), .B(n994), .Y(n993) );
  MXI2X1 U1919 ( .A(n995), .B(n953), .S0(n1883), .Y(n994) );
  MXI2X1 U1920 ( .A(n868), .B(n978), .S0(n1883), .Y(n992) );
  NAND2X1 U1921 ( .A(n996), .B(n997), .Y(addr_o[2]) );
  AOI221XL U1922 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N211 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N243 ), .B1(n865), .C0(n998), 
        .Y(n997) );
  OAI22X1 U1923 ( .A0(n999), .A1(n953), .B0(n1000), .B1(n951), .Y(n998) );
  AOI22X1 U1924 ( .A0(n919), .A1(n565), .B0(n878), .B1(\iexec_stage/BUS468[1] ), .Y(n1000) );
  AND2X1 U1925 ( .A(n1001), .B(n1002), .Y(n999) );
  AOI221XL U1926 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N178 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N114 ), .B1(n855), .C0(n1003), .Y(n996)
         );
  OAI2BB1X1 U1927 ( .A0N(n546), .A1N(n889), .B0(n1004), .Y(n1003) );
  MXI2X1 U1928 ( .A(n1005), .B(n1006), .S0(n585), .Y(n1004) );
  NOR2X1 U1929 ( .A(n861), .B(n546), .Y(n1006) );
  OAI2BB1X1 U1930 ( .A0N(n862), .A1N(n546), .B0(n863), .Y(n1005) );
  NAND4X1 U1931 ( .A(n1007), .B(n1008), .C(n1009), .D(n1010), .Y(addr_o[29])
         );
  AOI221XL U1932 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N205 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N141 ), .B1(n855), .C0(n1011), .Y(n1010) );
  OAI21X1 U1933 ( .A0(n1885), .A1(n988), .B0(n1012), .Y(n1011) );
  MXI2X1 U1934 ( .A(n1013), .B(n1014), .S0(n575), .Y(n1012) );
  NOR2X1 U1935 ( .A(n861), .B(n547), .Y(n1014) );
  NAND2X1 U1936 ( .A(n1015), .B(n863), .Y(n1013) );
  MXI2X1 U1937 ( .A(n862), .B(n868), .S0(n1885), .Y(n1015) );
  AOI22X1 U1938 ( .A0(n1016), .A1(n868), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N206 ), .B1(n871), .Y(n1009) );
  NAND2X1 U1939 ( .A(n973), .B(n986), .Y(n1008) );
  NAND4X1 U1940 ( .A(n1017), .B(n900), .C(n1018), .D(n882), .Y(n986) );
  NOR2X1 U1941 ( .A(n919), .B(n903), .Y(n1018) );
  AOI32X1 U1942 ( .A0(n878), .A1(n545), .A2(n1019), .B0(n990), .B1(n919), .Y(
        n1007) );
  CLKINVX1 U1943 ( .A(n1020), .Y(n1019) );
  NAND2X1 U1944 ( .A(n1021), .B(n1022), .Y(addr_o[28]) );
  AOI222XL U1945 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N204 ), .A1(n78), .B0(
        n868), .B1(n1023), .C0(n1024), .C1(n1025), .Y(n1022) );
  OAI221X1 U1946 ( .A0(n1026), .A1(n1027), .B0(n1028), .B1(n1029), .C0(n1030), 
        .Y(n1025) );
  NAND2X1 U1947 ( .A(\iexec_stage/MIPS_alu/mips_shifter/N205 ), .B(n1031), .Y(
        n1030) );
  NOR2X1 U1948 ( .A(n902), .B(n1032), .Y(n1028) );
  AOI31X1 U1949 ( .A0(n900), .A1(n881), .A2(n1017), .B0(n1033), .Y(n1032) );
  AOI222XL U1950 ( .A0(n879), .A1(n548), .B0(n919), .B1(n545), .C0(n878), .C1(
        n547), .Y(n1027) );
  OR2X1 U1951 ( .A(n1034), .B(n1035), .Y(n1023) );
  AOI221XL U1952 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N140 ), .A1(n855), .B0(
        n857), .B1(n548), .C0(n1036), .Y(n1021) );
  MXI2X1 U1953 ( .A(n1037), .B(n1038), .S0(n576), .Y(n1036) );
  NAND2X1 U1954 ( .A(n1886), .B(n978), .Y(n1038) );
  AOI21X1 U1955 ( .A0(n862), .A1(n548), .B0(n979), .Y(n1037) );
  NAND2X1 U1956 ( .A(n1039), .B(n1040), .Y(addr_o[27]) );
  AOI221XL U1957 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N204 ), .A1(n871), 
        .B0(\iexec_stage/MIPS_alu/mips_alu/N203 ), .B1(n78), .C0(n1041), .Y(
        n1040) );
  OAI22X1 U1958 ( .A0(n1042), .A1(n1043), .B0(n1044), .B1(n953), .Y(n1041) );
  NOR2X1 U1959 ( .A(n1045), .B(n1046), .Y(n1044) );
  AOI211X1 U1960 ( .A0(n903), .A1(n1047), .B0(n1048), .C0(n1049), .Y(n1042) );
  OAI22X1 U1961 ( .A0(n900), .A1(n1033), .B0(n1026), .B1(n1050), .Y(n1048) );
  AOI222XL U1962 ( .A0(n878), .A1(n548), .B0(n902), .B1(n545), .C0(n919), .C1(
        n547), .Y(n1050) );
  CLKINVX1 U1963 ( .A(n1051), .Y(n1026) );
  AOI221XL U1964 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N139 ), .A1(n855), .B0(
        n1052), .B1(n549), .C0(n1053), .Y(n1039) );
  MXI2X1 U1965 ( .A(n1054), .B(n1055), .S0(n577), .Y(n1053) );
  NAND2X1 U1966 ( .A(n1889), .B(n978), .Y(n1055) );
  AOI21X1 U1967 ( .A0(n862), .A1(n549), .B0(n979), .Y(n1054) );
  CLKINVX1 U1968 ( .A(n988), .Y(n1052) );
  AOI2BB1X1 U1969 ( .A0N(n980), .A1N(n1020), .B0(n857), .Y(n988) );
  NAND2X1 U1970 ( .A(n1056), .B(n1057), .Y(addr_o[26]) );
  AOI221XL U1971 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N203 ), .A1(n871), 
        .B0(\iexec_stage/MIPS_alu/mips_alu/N202 ), .B1(n78), .C0(n1058), .Y(
        n1057) );
  OAI22X1 U1972 ( .A0(n1059), .A1(n1043), .B0(n1060), .B1(n953), .Y(n1058) );
  AND2X1 U1973 ( .A(n1061), .B(n1062), .Y(n1060) );
  AOI221XL U1974 ( .A0(n1063), .A1(n1051), .B0(n873), .B1(n1047), .C0(n1049), 
        .Y(n1059) );
  CLKINVX1 U1975 ( .A(n1029), .Y(n1047) );
  NOR2BX1 U1976 ( .AN(n1033), .B(n1064), .Y(n1029) );
  OAI221X1 U1977 ( .A0(n1889), .A1(n905), .B0(n1891), .B1(n980), .C0(n1065), 
        .Y(n1063) );
  AOI222XL U1978 ( .A0(n919), .A1(n548), .B0(n902), .B1(n547), .C0(n903), .C1(
        n545), .Y(n1065) );
  AOI221XL U1979 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N138 ), .A1(n855), .B0(
        n857), .B1(n550), .C0(n1066), .Y(n1056) );
  MXI2X1 U1980 ( .A(n1067), .B(n1068), .S0(n578), .Y(n1066) );
  NAND2X1 U1981 ( .A(n1891), .B(n978), .Y(n1068) );
  AOI21X1 U1982 ( .A0(n862), .A1(n550), .B0(n979), .Y(n1067) );
  NAND2X1 U1983 ( .A(n1069), .B(n1070), .Y(addr_o[25]) );
  AOI221XL U1984 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N202 ), .A1(n871), 
        .B0(\iexec_stage/MIPS_alu/mips_alu/N201 ), .B1(n78), .C0(n1071), .Y(
        n1070) );
  OAI22X1 U1985 ( .A0(n1072), .A1(n1043), .B0(n1073), .B1(n953), .Y(n1071) );
  AND2X1 U1986 ( .A(n1074), .B(n1075), .Y(n1073) );
  AOI221XL U1987 ( .A0(n1076), .A1(n1051), .B0(n1064), .B1(n898), .C0(n1049), 
        .Y(n1072) );
  NOR2X1 U1988 ( .A(n1033), .B(n1017), .Y(n1049) );
  NOR2X1 U1989 ( .A(n1077), .B(n898), .Y(n1017) );
  NAND2X1 U1990 ( .A(n1078), .B(\iexec_stage/BUS468[31] ), .Y(n1033) );
  NOR2X1 U1991 ( .A(n1079), .B(n1881), .Y(n1064) );
  NAND2X1 U1992 ( .A(n1080), .B(n1081), .Y(n1076) );
  AOI222XL U1993 ( .A0(n903), .A1(n547), .B0(n873), .B1(n545), .C0(n902), .C1(
        n548), .Y(n1081) );
  AOI222XL U1994 ( .A0(n879), .A1(n551), .B0(n919), .B1(n549), .C0(n878), .C1(
        n550), .Y(n1080) );
  AOI221XL U1995 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N137 ), .A1(n855), .B0(
        n857), .B1(n551), .C0(n1082), .Y(n1069) );
  MXI2X1 U1996 ( .A(n1083), .B(n1084), .S0(n579), .Y(n1082) );
  NAND2X1 U1997 ( .A(n1892), .B(n978), .Y(n1084) );
  AOI21X1 U1998 ( .A0(n862), .A1(n551), .B0(n979), .Y(n1083) );
  NAND3X1 U1999 ( .A(n1085), .B(n1086), .C(n1087), .Y(addr_o[24]) );
  AOI221XL U2000 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N200 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N136 ), .B1(n855), .C0(n1088), .Y(n1087) );
  OAI2BB1X1 U2001 ( .A0N(n857), .A1N(n552), .B0(n1089), .Y(n1088) );
  MXI2X1 U2002 ( .A(n1090), .B(n1091), .S0(n580), .Y(n1089) );
  NOR2X1 U2003 ( .A(n861), .B(n552), .Y(n1091) );
  OAI2BB1X1 U2004 ( .A0N(n862), .A1N(n552), .B0(n863), .Y(n1090) );
  AOI222XL U2005 ( .A0(n990), .A1(n872), .B0(n1092), .B1(n1093), .C0(n868), 
        .C1(n1094), .Y(n1086) );
  NAND2X1 U2006 ( .A(n1095), .B(n1096), .Y(n1094) );
  NAND2X1 U2007 ( .A(n1097), .B(n1098), .Y(n1093) );
  AOI221XL U2008 ( .A0(n879), .A1(n552), .B0(n898), .B1(n545), .C0(n1099), .Y(
        n1098) );
  OAI22X1 U2009 ( .A0(n1892), .A1(n905), .B0(n1891), .B1(n883), .Y(n1099) );
  AOI222XL U2010 ( .A0(n903), .A1(n548), .B0(n873), .B1(n547), .C0(n902), .C1(
        n549), .Y(n1097) );
  AOI22X1 U2011 ( .A0(n973), .A1(n1077), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N201 ), .B1(n871), .Y(n1085) );
  OR2X1 U2012 ( .A(n1100), .B(n872), .Y(n1077) );
  NAND3X1 U2013 ( .A(n1101), .B(n1102), .C(n1103), .Y(addr_o[23]) );
  AOI221XL U2014 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N199 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N135 ), .B1(n855), .C0(n1104), .Y(n1103) );
  OAI2BB1X1 U2015 ( .A0N(n857), .A1N(n553), .B0(n1105), .Y(n1104) );
  MXI2X1 U2016 ( .A(n1106), .B(n1107), .S0(n581), .Y(n1105) );
  NOR2X1 U2017 ( .A(n861), .B(n553), .Y(n1107) );
  OAI2BB1X1 U2018 ( .A0N(n862), .A1N(n553), .B0(n863), .Y(n1106) );
  AOI222XL U2019 ( .A0(n990), .A1(n897), .B0(n1092), .B1(n1108), .C0(n868), 
        .C1(n1109), .Y(n1102) );
  OR2X1 U2020 ( .A(n1110), .B(n1111), .Y(n1109) );
  NAND2X1 U2021 ( .A(n1112), .B(n1113), .Y(n1108) );
  AOI221XL U2022 ( .A0(n898), .A1(n547), .B0(n872), .B1(n545), .C0(n1114), .Y(
        n1113) );
  OAI22X1 U2023 ( .A0(n1889), .A1(n881), .B0(n1886), .B1(n900), .Y(n1114) );
  AOI221XL U2024 ( .A0(n878), .A1(n552), .B0(n879), .B1(n553), .C0(n1115), .Y(
        n1112) );
  OAI22X1 U2025 ( .A0(n1892), .A1(n883), .B0(n1891), .B1(n882), .Y(n1115) );
  AOI22X1 U2026 ( .A0(n973), .A1(n1100), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N200 ), .B1(n871), .Y(n1101) );
  OR2X1 U2027 ( .A(n1116), .B(n897), .Y(n1100) );
  NAND3X1 U2028 ( .A(n1117), .B(n1118), .C(n1119), .Y(addr_o[22]) );
  AOI221XL U2029 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N198 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N134 ), .B1(n855), .C0(n1120), .Y(n1119) );
  OAI2BB1X1 U2030 ( .A0N(n857), .A1N(n554), .B0(n1121), .Y(n1120) );
  MXI2X1 U2031 ( .A(n1122), .B(n1123), .S0(n582), .Y(n1121) );
  NOR2X1 U2032 ( .A(n861), .B(n554), .Y(n1123) );
  OAI2BB1X1 U2033 ( .A0N(n862), .A1N(n554), .B0(n863), .Y(n1122) );
  AOI221XL U2034 ( .A0(n990), .A1(n1124), .B0(n868), .B1(n1125), .C0(n1126), 
        .Y(n1118) );
  AOI31X1 U2035 ( .A0(n1127), .A1(n1128), .A2(n1129), .B0(n1130), .Y(n1126) );
  AOI221XL U2036 ( .A0(n878), .A1(n553), .B0(n879), .B1(n554), .C0(n1131), .Y(
        n1129) );
  OAI22X1 U2037 ( .A0(n1893), .A1(n883), .B0(n1892), .B1(n882), .Y(n1131) );
  AOI222XL U2038 ( .A0(n872), .A1(n547), .B0(n897), .B1(n545), .C0(n898), .C1(
        n548), .Y(n1128) );
  AOI22X1 U2039 ( .A0(n873), .A1(n549), .B0(n903), .B1(n550), .Y(n1127) );
  OR2X1 U2040 ( .A(n1132), .B(n1133), .Y(n1125) );
  AOI22X1 U2041 ( .A0(n973), .A1(n1116), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N199 ), .B1(n871), .Y(n1117) );
  OR2X1 U2042 ( .A(n1134), .B(n1124), .Y(n1116) );
  NAND3X1 U2043 ( .A(n1135), .B(n1136), .C(n1137), .Y(addr_o[21]) );
  AOI221XL U2044 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N197 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N133 ), .B1(n855), .C0(n1138), .Y(n1137) );
  OAI2BB1X1 U2045 ( .A0N(n857), .A1N(n555), .B0(n1139), .Y(n1138) );
  MXI2X1 U2046 ( .A(n1140), .B(n1141), .S0(n583), .Y(n1139) );
  NOR2X1 U2047 ( .A(n861), .B(n555), .Y(n1141) );
  OAI2BB1X1 U2048 ( .A0N(n862), .A1N(n555), .B0(n863), .Y(n1140) );
  AOI222XL U2049 ( .A0(n1142), .A1(n990), .B0(n1092), .B1(n1143), .C0(n868), 
        .C1(n1144), .Y(n1136) );
  OR2X1 U2050 ( .A(n1145), .B(n1146), .Y(n1144) );
  NAND4X1 U2051 ( .A(n1147), .B(n1148), .C(n1149), .D(n1150), .Y(n1143) );
  AOI222XL U2052 ( .A0(n898), .A1(n549), .B0(n1124), .B1(n545), .C0(n897), 
        .C1(n547), .Y(n1150) );
  AOI22X1 U2053 ( .A0(n872), .A1(n548), .B0(n873), .B1(n550), .Y(n1149) );
  AOI222XL U2054 ( .A0(n919), .A1(n553), .B0(n902), .B1(n552), .C0(n903), .C1(
        n551), .Y(n1148) );
  AOI22X1 U2055 ( .A0(n878), .A1(n554), .B0(n879), .B1(n555), .Y(n1147) );
  AOI22X1 U2056 ( .A0(n973), .A1(n1134), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N198 ), .B1(n871), .Y(n1135) );
  OR2X1 U2057 ( .A(n1151), .B(n1142), .Y(n1134) );
  NAND3X1 U2058 ( .A(n1152), .B(n1153), .C(n1154), .Y(addr_o[20]) );
  AOI221XL U2059 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N196 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N132 ), .B1(n855), .C0(n1155), .Y(n1154) );
  OAI21X1 U2060 ( .A0(n1898), .A1(n982), .B0(n1156), .Y(n1155) );
  MXI2X1 U2061 ( .A(n1157), .B(n1158), .S0(n584), .Y(n1156) );
  NOR2X1 U2062 ( .A(n861), .B(n556), .Y(n1158) );
  OAI2BB1X1 U2063 ( .A0N(n862), .A1N(n556), .B0(n863), .Y(n1157) );
  AOI222XL U2064 ( .A0(n1159), .A1(n1092), .B0(n868), .B1(n1160), .C0(n1161), 
        .C1(n990), .Y(n1153) );
  NAND2X1 U2065 ( .A(n1162), .B(n1163), .Y(n1160) );
  NAND4X1 U2066 ( .A(n1164), .B(n1165), .C(n1166), .D(n1167), .Y(n1159) );
  AOI222XL U2067 ( .A0(n897), .A1(n548), .B0(n1124), .B1(n547), .C0(n1142), 
        .C1(n545), .Y(n1167) );
  AOI222XL U2068 ( .A0(n873), .A1(n551), .B0(n898), .B1(n550), .C0(n872), .C1(
        n549), .Y(n1166) );
  AOI222XL U2069 ( .A0(n919), .A1(n554), .B0(n902), .B1(n553), .C0(n903), .C1(
        n552), .Y(n1165) );
  AOI22X1 U2070 ( .A0(n878), .A1(n555), .B0(n879), .B1(n556), .Y(n1164) );
  AOI22X1 U2071 ( .A0(n973), .A1(n1151), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N197 ), .B1(n871), .Y(n1152) );
  NAND3BX1 U2072 ( .AN(n1168), .B(n1169), .C(n1170), .Y(n1151) );
  NAND2X1 U2073 ( .A(n1171), .B(n1172), .Y(addr_o[1]) );
  AOI221XL U2074 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N210 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N242 ), .B1(n865), .C0(n1173), 
        .Y(n1172) );
  OAI32X1 U2075 ( .A0(n951), .A1(n1927), .A2(n905), .B0(n1926), .B1(n967), .Y(
        n1173) );
  AOI221XL U2076 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N177 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N113 ), .B1(n855), .C0(n1174), .Y(n1171) );
  MXI2X1 U2077 ( .A(n1175), .B(n1176), .S0(n596), .Y(n1174) );
  MXI2X1 U2078 ( .A(n868), .B(n978), .S0(n1926), .Y(n1176) );
  NOR2X1 U2079 ( .A(n979), .B(n1177), .Y(n1175) );
  MXI2X1 U2080 ( .A(n995), .B(n953), .S0(n1926), .Y(n1177) );
  NAND3X1 U2081 ( .A(n1178), .B(n1179), .C(n1180), .Y(addr_o[19]) );
  AOI221XL U2082 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N195 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N131 ), .B1(n855), .C0(n1181), .Y(n1180) );
  OAI21X1 U2083 ( .A0(n1899), .A1(n982), .B0(n1182), .Y(n1181) );
  MXI2X1 U2084 ( .A(n1183), .B(n1184), .S0(n586), .Y(n1182) );
  NOR2X1 U2085 ( .A(n861), .B(n557), .Y(n1184) );
  OAI2BB1X1 U2086 ( .A0N(n862), .A1N(n557), .B0(n863), .Y(n1183) );
  AOI222XL U2087 ( .A0(n973), .A1(n1168), .B0(n868), .B1(n1185), .C0(n1186), 
        .C1(n1187), .Y(n1179) );
  NAND2X1 U2088 ( .A(n1188), .B(n1189), .Y(n1185) );
  OR2X1 U2089 ( .A(n1190), .B(n1191), .Y(n1168) );
  AOI22X1 U2090 ( .A0(n1192), .A1(n1092), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N196 ), .B1(n871), .Y(n1178) );
  NAND4X1 U2091 ( .A(n1193), .B(n1194), .C(n1195), .D(n1196), .Y(n1192) );
  AOI222XL U2092 ( .A0(n1142), .A1(n547), .B0(n1161), .B1(n545), .C0(n1124), 
        .C1(n548), .Y(n1196) );
  AOI222XL U2093 ( .A0(n872), .A1(n550), .B0(n897), .B1(n549), .C0(n898), .C1(
        n551), .Y(n1195) );
  AOI222XL U2094 ( .A0(n903), .A1(n553), .B0(n873), .B1(n552), .C0(n902), .C1(
        n554), .Y(n1194) );
  AOI222XL U2095 ( .A0(n879), .A1(n557), .B0(n919), .B1(n555), .C0(n878), .C1(
        n556), .Y(n1193) );
  NAND3X1 U2096 ( .A(n1197), .B(n1198), .C(n1199), .Y(addr_o[18]) );
  AOI221XL U2097 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N194 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N130 ), .B1(n855), .C0(n1200), .Y(n1199) );
  OAI21X1 U2098 ( .A0(n1901), .A1(n982), .B0(n1201), .Y(n1200) );
  MXI2X1 U2099 ( .A(n1202), .B(n1203), .S0(n587), .Y(n1201) );
  NOR2X1 U2100 ( .A(n861), .B(n558), .Y(n1203) );
  OAI2BB1X1 U2101 ( .A0N(n862), .A1N(n558), .B0(n863), .Y(n1202) );
  AOI222XL U2102 ( .A0(n973), .A1(n1190), .B0(n868), .B1(n1204), .C0(n1191), 
        .C1(n1186), .Y(n1198) );
  NAND2X1 U2103 ( .A(n1205), .B(n1206), .Y(n1204) );
  AOI22X1 U2104 ( .A0(n1207), .A1(n1092), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N195 ), .B1(n871), .Y(n1197) );
  NAND4X1 U2105 ( .A(n1208), .B(n1209), .C(n1210), .D(n1211), .Y(n1207) );
  AOI221XL U2106 ( .A0(n1187), .A1(n545), .B0(n1161), .B1(n547), .C0(n1212), 
        .Y(n1211) );
  OAI22X1 U2107 ( .A0(n1886), .A1(n1213), .B0(n1889), .B1(n876), .Y(n1212) );
  AOI222XL U2108 ( .A0(n872), .A1(n551), .B0(n897), .B1(n550), .C0(n898), .C1(
        n552), .Y(n1210) );
  AOI222XL U2109 ( .A0(n903), .A1(n554), .B0(n873), .B1(n553), .C0(n902), .C1(
        n555), .Y(n1209) );
  AOI222XL U2110 ( .A0(n879), .A1(n558), .B0(n919), .B1(n556), .C0(n878), .C1(
        n557), .Y(n1208) );
  NAND3X1 U2111 ( .A(n1214), .B(n1215), .C(n1216), .Y(addr_o[17]) );
  AOI221XL U2112 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N193 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N129 ), .B1(n855), .C0(n1217), .Y(n1216) );
  OAI21X1 U2113 ( .A0(n1903), .A1(n982), .B0(n1218), .Y(n1217) );
  MXI2X1 U2114 ( .A(n1219), .B(n1220), .S0(n588), .Y(n1218) );
  NOR2X1 U2115 ( .A(n861), .B(n559), .Y(n1220) );
  OAI2BB1X1 U2116 ( .A0N(n862), .A1N(n559), .B0(n863), .Y(n1219) );
  AOI222XL U2117 ( .A0(n973), .A1(n1190), .B0(n868), .B1(n1221), .C0(n1222), 
        .C1(n990), .Y(n1215) );
  NOR2X1 U2118 ( .A(n981), .B(n1881), .Y(n990) );
  OR2X1 U2119 ( .A(n1223), .B(n1224), .Y(n1221) );
  AOI22X1 U2120 ( .A0(n1226), .A1(n1092), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N194 ), .B1(n871), .Y(n1214) );
  NAND4X1 U2121 ( .A(n1227), .B(n1228), .C(n1229), .D(n1230), .Y(n1226) );
  AOI221XL U2122 ( .A0(n1191), .A1(n545), .B0(n1187), .B1(n547), .C0(n1231), 
        .Y(n1230) );
  OAI22X1 U2123 ( .A0(n1891), .A1(n876), .B0(n1886), .B1(n1170), .Y(n1231) );
  AOI222XL U2124 ( .A0(n898), .A1(n553), .B0(n1142), .B1(n549), .C0(n897), 
        .C1(n551), .Y(n1229) );
  AOI221XL U2125 ( .A0(n872), .A1(n552), .B0(n873), .B1(n554), .C0(n1232), .Y(
        n1228) );
  OAI22X1 U2126 ( .A0(n1897), .A1(n881), .B0(n1898), .B1(n882), .Y(n1232) );
  AOI222XL U2127 ( .A0(n879), .A1(n559), .B0(n919), .B1(n557), .C0(n878), .C1(
        n558), .Y(n1227) );
  NAND3X1 U2128 ( .A(n1233), .B(n1234), .C(n1235), .Y(addr_o[16]) );
  AOI221XL U2129 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N192 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N128 ), .B1(n855), .C0(n1236), .Y(n1235) );
  OAI21X1 U2130 ( .A0(n1906), .A1(n982), .B0(n1237), .Y(n1236) );
  MXI2X1 U2131 ( .A(n1238), .B(n1239), .S0(n589), .Y(n1237) );
  NOR2X1 U2132 ( .A(n861), .B(n567), .Y(n1239) );
  OAI2BB1X1 U2133 ( .A0N(n862), .A1N(n567), .B0(n863), .Y(n1238) );
  AOI222XL U2134 ( .A0(n973), .A1(\iexec_stage/BUS476[4] ), .B0(n868), .B1(
        n1240), .C0(n1225), .C1(n1186), .Y(n1234) );
  NOR2X1 U2135 ( .A(n1130), .B(n1881), .Y(n1186) );
  CLKINVX1 U2136 ( .A(n1092), .Y(n1130) );
  OR2X1 U2137 ( .A(n1241), .B(n1242), .Y(n1240) );
  NOR2X1 U2138 ( .A(n1243), .B(n1881), .Y(n973) );
  AOI22X1 U2139 ( .A0(n1244), .A1(n1092), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N193 ), .B1(n871), .Y(n1233) );
  NAND2X1 U2140 ( .A(n1243), .B(n981), .Y(n1092) );
  CLKINVX1 U2141 ( .A(n864), .Y(n981) );
  NAND4X1 U2142 ( .A(n1245), .B(n1246), .C(n1247), .D(n1248), .Y(n1244) );
  AOI221XL U2143 ( .A0(n1222), .A1(n545), .B0(n1191), .B1(n547), .C0(n1249), 
        .Y(n1248) );
  OAI22X1 U2144 ( .A0(n1889), .A1(n1170), .B0(n1886), .B1(n1169), .Y(n1249) );
  AOI221XL U2145 ( .A0(n1124), .A1(n551), .B0(n1142), .B1(n550), .C0(n1250), 
        .Y(n1247) );
  OAI22X1 U2146 ( .A0(n1896), .A1(n877), .B0(n1893), .B1(n875), .Y(n1250) );
  AOI221XL U2147 ( .A0(n872), .A1(n553), .B0(n873), .B1(n555), .C0(n1251), .Y(
        n1246) );
  OAI22X1 U2148 ( .A0(n1898), .A1(n881), .B0(n1899), .B1(n882), .Y(n1251) );
  AOI222XL U2149 ( .A0(n879), .A1(n567), .B0(n919), .B1(n558), .C0(n878), .C1(
        n559), .Y(n1245) );
  NAND4X1 U2150 ( .A(n1252), .B(n1253), .C(n1254), .D(n1255), .Y(addr_o[15])
         );
  AOI221XL U2151 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N191 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N127 ), .B1(n855), .C0(n1256), .Y(n1255) );
  OAI21X1 U2152 ( .A0(n1909), .A1(n982), .B0(n1257), .Y(n1256) );
  MXI2X1 U2153 ( .A(n1258), .B(n1259), .S0(n590), .Y(n1257) );
  NOR2X1 U2154 ( .A(\iexec_stage/BUS468[15] ), .B(n861), .Y(n1259) );
  OAI2BB1X1 U2155 ( .A0N(n862), .A1N(\iexec_stage/BUS468[15] ), .B0(n863), .Y(
        n1258) );
  AOI22X1 U2156 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N224 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N256 ), .B1(n865), .Y(n1254) );
  OAI21X1 U2157 ( .A0(n1260), .A1(n1261), .B0(n868), .Y(n1253) );
  NAND2X1 U2158 ( .A(n871), .B(n1262), .Y(n1252) );
  NAND4X1 U2159 ( .A(n1263), .B(n1264), .C(n1265), .D(n1266), .Y(n1262) );
  AOI221XL U2160 ( .A0(n1225), .A1(n565), .B0(n1222), .B1(
        \iexec_stage/BUS468[1] ), .C0(n1267), .Y(n1266) );
  OAI22X1 U2161 ( .A0(n1924), .A1(n1169), .B0(n1925), .B1(n1268), .Y(n1267) );
  AND2X1 U2162 ( .A(n1269), .B(n1270), .Y(n1225) );
  AOI221XL U2163 ( .A0(n1161), .A1(n543), .B0(n1124), .B1(n541), .C0(n1271), 
        .Y(n1265) );
  OAI22X1 U2164 ( .A0(n1919), .A1(n875), .B0(n1921), .B1(n1213), .Y(n1271) );
  AOI221XL U2165 ( .A0(n898), .A1(\iexec_stage/BUS468[9] ), .B0(n872), .B1(
        n539), .C0(n1272), .Y(n1264) );
  OAI22X1 U2166 ( .A0(n1913), .A1(n882), .B0(n1916), .B1(n900), .Y(n1272) );
  AOI221XL U2167 ( .A0(n903), .A1(n563), .B0(n919), .B1(n561), .C0(n1273), .Y(
        n1263) );
  OAI22X1 U2168 ( .A0(n1909), .A1(n980), .B0(n1911), .B1(n905), .Y(n1273) );
  NAND4X1 U2169 ( .A(n1274), .B(n1275), .C(n1276), .D(n1277), .Y(addr_o[14])
         );
  AOI221XL U2170 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N190 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N126 ), .B1(n855), .C0(n1278), .Y(n1277) );
  OAI21X1 U2171 ( .A0(n1911), .A1(n982), .B0(n1279), .Y(n1278) );
  MXI2X1 U2172 ( .A(n1280), .B(n1281), .S0(n591), .Y(n1279) );
  NOR2X1 U2173 ( .A(n861), .B(n560), .Y(n1281) );
  OAI2BB1X1 U2174 ( .A0N(n862), .A1N(n560), .B0(n863), .Y(n1280) );
  AOI22X1 U2175 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N223 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N255 ), .B1(n865), .Y(n1276) );
  OAI2BB1X1 U2176 ( .A0N(n1282), .A1N(n1283), .B0(n868), .Y(n1275) );
  NAND2X1 U2177 ( .A(n871), .B(n1284), .Y(n1274) );
  NAND4X1 U2178 ( .A(n1285), .B(n1286), .C(n1287), .D(n1288), .Y(n1284) );
  AOI221XL U2179 ( .A0(n1222), .A1(n565), .B0(n1191), .B1(
        \iexec_stage/BUS468[1] ), .C0(n1289), .Y(n1288) );
  OAI22X1 U2180 ( .A0(n1924), .A1(n1170), .B0(n1925), .B1(n1169), .Y(n1289) );
  AND2X1 U2181 ( .A(n1269), .B(n1290), .Y(n1222) );
  AOI221XL U2182 ( .A0(n1124), .A1(n542), .B0(n1142), .B1(n543), .C0(n1291), 
        .Y(n1287) );
  OAI22X1 U2183 ( .A0(n1918), .A1(n877), .B0(n1920), .B1(n875), .Y(n1291) );
  AOI221XL U2184 ( .A0(n872), .A1(n540), .B0(n873), .B1(
        \iexec_stage/BUS468[9] ), .C0(n1292), .Y(n1286) );
  OAI22X1 U2185 ( .A0(n1916), .A1(n881), .B0(n1915), .B1(n882), .Y(n1292) );
  AOI222XL U2186 ( .A0(n879), .A1(n560), .B0(n919), .B1(n562), .C0(n878), .C1(
        n561), .Y(n1285) );
  NAND4X1 U2187 ( .A(n1293), .B(n1294), .C(n1295), .D(n1296), .Y(addr_o[13])
         );
  AOI221XL U2188 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N189 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N125 ), .B1(n855), .C0(n1297), .Y(n1296) );
  OAI21X1 U2189 ( .A0(n1912), .A1(n982), .B0(n1298), .Y(n1297) );
  MXI2X1 U2190 ( .A(n1299), .B(n1300), .S0(n592), .Y(n1298) );
  NOR2X1 U2191 ( .A(n861), .B(n561), .Y(n1300) );
  OAI2BB1X1 U2192 ( .A0N(n862), .A1N(n561), .B0(n863), .Y(n1299) );
  AOI22X1 U2193 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N222 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N254 ), .B1(n865), .Y(n1295) );
  OAI2BB1X1 U2194 ( .A0N(n1301), .A1N(n1302), .B0(n868), .Y(n1294) );
  NAND2X1 U2195 ( .A(n871), .B(n1303), .Y(n1293) );
  NAND4X1 U2196 ( .A(n1304), .B(n1305), .C(n1306), .D(n1307), .Y(n1303) );
  AOI221XL U2197 ( .A0(n1191), .A1(n565), .B0(n1187), .B1(
        \iexec_stage/BUS468[1] ), .C0(n1308), .Y(n1307) );
  OAI22X1 U2198 ( .A0(n1922), .A1(n876), .B0(n1925), .B1(n1170), .Y(n1308) );
  CLKINVX1 U2199 ( .A(n1268), .Y(n1191) );
  NAND2X1 U2200 ( .A(n1270), .B(n1309), .Y(n1268) );
  AOI222XL U2201 ( .A0(n898), .A1(n540), .B0(n1142), .B1(n544), .C0(n897), 
        .C1(n542), .Y(n1306) );
  AOI221XL U2202 ( .A0(n872), .A1(n541), .B0(n873), .B1(n539), .C0(n1310), .Y(
        n1305) );
  OAI22X1 U2203 ( .A0(n1917), .A1(n881), .B0(n1916), .B1(n882), .Y(n1310) );
  AOI222XL U2204 ( .A0(n879), .A1(n561), .B0(n919), .B1(n563), .C0(n878), .C1(
        n562), .Y(n1304) );
  NAND4X1 U2205 ( .A(n1311), .B(n1312), .C(n1313), .D(n1314), .Y(addr_o[12])
         );
  AOI221XL U2206 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N188 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N124 ), .B1(n855), .C0(n1315), .Y(n1314) );
  OAI21X1 U2207 ( .A0(n1913), .A1(n982), .B0(n1316), .Y(n1315) );
  MXI2X1 U2208 ( .A(n1317), .B(n1318), .S0(n593), .Y(n1316) );
  NOR2X1 U2209 ( .A(n861), .B(n562), .Y(n1318) );
  OAI2BB1X1 U2210 ( .A0N(n862), .A1N(n562), .B0(n863), .Y(n1317) );
  AOI22X1 U2211 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N221 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N253 ), .B1(n865), .Y(n1313) );
  OAI2BB1X1 U2212 ( .A0N(n1319), .A1N(n1320), .B0(n868), .Y(n1312) );
  NAND2X1 U2213 ( .A(n871), .B(n1321), .Y(n1311) );
  NAND4X1 U2214 ( .A(n1322), .B(n1323), .C(n1324), .D(n1325), .Y(n1321) );
  AOI221XL U2215 ( .A0(n1187), .A1(n565), .B0(n1161), .B1(
        \iexec_stage/BUS468[1] ), .C0(n1326), .Y(n1325) );
  OAI22X1 U2216 ( .A0(n1925), .A1(n1213), .B0(n1924), .B1(n876), .Y(n1326) );
  CLKINVX1 U2217 ( .A(n1169), .Y(n1187) );
  NAND2X1 U2218 ( .A(n1290), .B(n1309), .Y(n1169) );
  AOI222XL U2219 ( .A0(n872), .A1(n542), .B0(n897), .B1(n543), .C0(n898), .C1(
        n541), .Y(n1324) );
  AOI222XL U2220 ( .A0(n903), .A1(n539), .B0(n873), .B1(n540), .C0(n902), .C1(
        \iexec_stage/BUS468[9] ), .Y(n1323) );
  AOI222XL U2221 ( .A0(n879), .A1(n562), .B0(n919), .B1(n564), .C0(n878), .C1(
        n563), .Y(n1322) );
  NAND4X1 U2222 ( .A(n1327), .B(n1328), .C(n1329), .D(n1330), .Y(addr_o[11])
         );
  AOI221XL U2223 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N187 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N123 ), .B1(n855), .C0(n1331), .Y(n1330) );
  OAI21X1 U2224 ( .A0(n1915), .A1(n982), .B0(n1332), .Y(n1331) );
  MXI2X1 U2225 ( .A(n1333), .B(n1334), .S0(n594), .Y(n1332) );
  NOR2X1 U2226 ( .A(n861), .B(n563), .Y(n1334) );
  OAI2BB1X1 U2227 ( .A0N(n862), .A1N(n563), .B0(n863), .Y(n1333) );
  AOI22X1 U2228 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N220 ), .A1(n864), 
        .B0(\iexec_stage/MIPS_alu/mips_shifter/N252 ), .B1(n865), .Y(n1329) );
  OAI21X1 U2229 ( .A0(n1335), .A1(n1336), .B0(n868), .Y(n1328) );
  NAND2X1 U2230 ( .A(n871), .B(n1337), .Y(n1327) );
  NAND4X1 U2231 ( .A(n1338), .B(n1339), .C(n1340), .D(n1341), .Y(n1337) );
  AOI222XL U2232 ( .A0(n1142), .A1(\iexec_stage/BUS468[1] ), .B0(n1161), .B1(
        n565), .C0(n1124), .C1(n546), .Y(n1341) );
  CLKINVX1 U2233 ( .A(n1170), .Y(n1161) );
  NAND2X1 U2234 ( .A(n1269), .B(n1342), .Y(n1170) );
  AOI222XL U2235 ( .A0(n872), .A1(n543), .B0(n897), .B1(n544), .C0(n898), .C1(
        n542), .Y(n1340) );
  AOI222XL U2236 ( .A0(n903), .A1(n540), .B0(n873), .B1(n541), .C0(n902), .C1(
        n539), .Y(n1339) );
  AOI222XL U2237 ( .A0(n879), .A1(n563), .B0(n919), .B1(
        \iexec_stage/BUS468[9] ), .C0(n878), .C1(n564), .Y(n1338) );
  NAND3X1 U2238 ( .A(n1343), .B(n1344), .C(n1345), .Y(addr_o[10]) );
  AOI221XL U2239 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N186 ), .A1(n78), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N122 ), .B1(n855), .C0(n1346), .Y(n1345) );
  OAI2BB1X1 U2240 ( .A0N(n857), .A1N(n564), .B0(n1347), .Y(n1346) );
  MXI2X1 U2241 ( .A(n1348), .B(n1349), .S0(n595), .Y(n1347) );
  NOR2X1 U2242 ( .A(n861), .B(n564), .Y(n1349) );
  CLKINVX1 U2243 ( .A(n978), .Y(n861) );
  OAI2BB1X1 U2244 ( .A0N(n862), .A1N(n564), .B0(n863), .Y(n1348) );
  AOI22X1 U2245 ( .A0(n868), .A1(n1350), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/N219 ), .B1(n864), .Y(n1344) );
  NOR2X1 U2246 ( .A(n1079), .B(n1043), .Y(n864) );
  OR2X1 U2247 ( .A(n1351), .B(n1352), .Y(n1350) );
  AOI22X1 U2248 ( .A0(\iexec_stage/MIPS_alu/mips_shifter/N251 ), .A1(n865), 
        .B0(n871), .B1(n1353), .Y(n1343) );
  NAND4X1 U2249 ( .A(n1354), .B(n1355), .C(n1356), .D(n1357), .Y(n1353) );
  AOI222XL U2250 ( .A0(n897), .A1(n546), .B0(n1124), .B1(
        \iexec_stage/BUS468[1] ), .C0(n1142), .C1(n565), .Y(n1357) );
  CLKINVX1 U2251 ( .A(n1213), .Y(n1142) );
  NAND2X1 U2252 ( .A(n1269), .B(n1358), .Y(n1213) );
  NOR2X1 U2253 ( .A(n574), .B(n596), .Y(n1269) );
  CLKINVX1 U2254 ( .A(n876), .Y(n1124) );
  NAND2X1 U2255 ( .A(n1309), .B(n1342), .Y(n876) );
  CLKINVX1 U2256 ( .A(n875), .Y(n897) );
  NAND2X1 U2257 ( .A(n1309), .B(n1358), .Y(n875) );
  NOR2X1 U2258 ( .A(n574), .B(\iexec_stage/BUS476[1] ), .Y(n1309) );
  AOI222XL U2259 ( .A0(n873), .A1(n542), .B0(n898), .B1(n543), .C0(n872), .C1(
        n544), .Y(n1356) );
  CLKINVX1 U2260 ( .A(n901), .Y(n872) );
  NAND2X1 U2261 ( .A(n1270), .B(n1359), .Y(n901) );
  CLKINVX1 U2262 ( .A(n877), .Y(n898) );
  NAND2X1 U2263 ( .A(n1359), .B(n1290), .Y(n877) );
  CLKINVX1 U2264 ( .A(n900), .Y(n873) );
  NAND2X1 U2265 ( .A(n1270), .B(n1360), .Y(n900) );
  AND2X1 U2266 ( .A(n1361), .B(\iexec_stage/BUS476[2] ), .Y(n1270) );
  AOI222XL U2267 ( .A0(n919), .A1(n539), .B0(n902), .B1(n540), .C0(n903), .C1(
        n541), .Y(n1355) );
  CLKINVX1 U2268 ( .A(n881), .Y(n903) );
  NAND2X1 U2269 ( .A(n1290), .B(n1360), .Y(n881) );
  AND2X1 U2270 ( .A(n1362), .B(\iexec_stage/BUS476[2] ), .Y(n1290) );
  CLKINVX1 U2271 ( .A(n882), .Y(n902) );
  NAND2X1 U2272 ( .A(n1359), .B(n1342), .Y(n882) );
  CLKINVX1 U2273 ( .A(n883), .Y(n919) );
  NAND2X1 U2274 ( .A(n1359), .B(n1358), .Y(n883) );
  NOR2X1 U2275 ( .A(n596), .B(\iexec_stage/BUS476[3] ), .Y(n1359) );
  AOI22X1 U2276 ( .A0(n878), .A1(\iexec_stage/BUS468[9] ), .B0(n879), .B1(n564), .Y(n1354) );
  CLKINVX1 U2277 ( .A(n980), .Y(n879) );
  CLKINVX1 U2278 ( .A(n905), .Y(n878) );
  NAND2X1 U2279 ( .A(n1360), .B(n1342), .Y(n905) );
  AND2X1 U2280 ( .A(n1361), .B(n585), .Y(n1342) );
  NOR2X1 U2281 ( .A(n597), .B(\iexec_stage/BUS476[4] ), .Y(n1361) );
  CLKINVX1 U2282 ( .A(n951), .Y(n871) );
  CLKINVX1 U2283 ( .A(n1243), .Y(n865) );
  NAND2X1 U2284 ( .A(n1078), .B(n1024), .Y(n1243) );
  NAND2X1 U2285 ( .A(n1363), .B(n1364), .Y(addr_o[0]) );
  AOI221XL U2286 ( .A0(n889), .A1(n565), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N176 ), .B1(n78), .C0(n1365), .Y(n1364)
         );
  OAI32X1 U2287 ( .A0(n1366), .A1(n1367), .A2(n1368), .B0(
        \iexec_stage/MIPS_alu/mips_shifter/n511 ), .B1(n1020), .Y(n1365) );
  NAND2X1 U2288 ( .A(n1024), .B(n1051), .Y(n1020) );
  NAND2X1 U2289 ( .A(n1079), .B(n1369), .Y(n1051) );
  NAND3X1 U2290 ( .A(n288), .B(n40), .C(n287), .Y(n1079) );
  AOI2BB1X1 U2291 ( .A0N(\iexec_stage/BUS476[31] ), .A1N(n1881), .B0(n1370), 
        .Y(n1367) );
  AOI222XL U2292 ( .A0(\iexec_stage/BUS476[31] ), .A1(n1881), .B0(n1371), .B1(
        \iexec_stage/BUS476[30] ), .C0(n1883), .C1(n1372), .Y(n1370) );
  NAND2X1 U2293 ( .A(n1373), .B(n1374), .Y(\iexec_stage/BUS476[30] ) );
  AOI222XL U2294 ( .A0(cop_addr_o[30]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[30]), .C0(BUS7101[30]), .C1(n1377), .Y(n1374) );
  AOI222XL U2295 ( .A0(\iexec_stage/BUS2332[30] ), .A1(n1378), .B0(BUS7231[30]), .B1(n1379), .C0(n1380), .C1(n71), .Y(n1373) );
  OR2X1 U2296 ( .A(n1372), .B(n1883), .Y(n1371) );
  CLKINVX1 U2297 ( .A(n545), .Y(n1883) );
  OAI221X1 U2298 ( .A0(n1381), .A1(n1382), .B0(n1383), .B1(n1384), .C0(n1385), 
        .Y(n545) );
  AOI22X1 U2299 ( .A0(cop_addr_o[30]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[30]), .Y(n1385) );
  CLKINVX1 U2300 ( .A(BUS7231[30]), .Y(n1382) );
  OAI32X1 U2301 ( .A0(n1035), .A1(n1388), .A2(n1016), .B0(n575), .B1(n547), 
        .Y(n1372) );
  CLKINVX1 U2302 ( .A(\iexec_stage/BUS476[29] ), .Y(n575) );
  NOR2X1 U2303 ( .A(n1885), .B(\iexec_stage/BUS476[29] ), .Y(n1016) );
  NAND2X1 U2304 ( .A(n1389), .B(n1390), .Y(\iexec_stage/BUS476[29] ) );
  AOI222XL U2305 ( .A0(cop_addr_o[29]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[29]), .C0(BUS7101[29]), .C1(n1377), .Y(n1390) );
  AOI222XL U2306 ( .A0(\iexec_stage/BUS2332[29] ), .A1(n1378), .B0(BUS7231[29]), .B1(n1379), .C0(n1380), .C1(n72), .Y(n1389) );
  CLKINVX1 U2307 ( .A(n547), .Y(n1885) );
  OAI221X1 U2308 ( .A0(n1381), .A1(n1391), .B0(n1383), .B1(n1392), .C0(n1393), 
        .Y(n547) );
  AOI22X1 U2309 ( .A0(cop_addr_o[29]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[29]), .Y(n1393) );
  CLKINVX1 U2310 ( .A(BUS7231[29]), .Y(n1391) );
  AOI211X1 U2311 ( .A0(n1394), .A1(n1061), .B0(n1045), .C0(n1034), .Y(n1388)
         );
  NOR2X1 U2312 ( .A(n548), .B(n576), .Y(n1034) );
  CLKINVX1 U2313 ( .A(\iexec_stage/BUS476[28] ), .Y(n576) );
  NOR2X1 U2314 ( .A(n549), .B(n577), .Y(n1045) );
  CLKINVX1 U2315 ( .A(\iexec_stage/BUS476[27] ), .Y(n577) );
  NAND2X1 U2316 ( .A(n550), .B(n578), .Y(n1061) );
  CLKINVX1 U2317 ( .A(\iexec_stage/BUS476[26] ), .Y(n578) );
  AOI31X1 U2318 ( .A0(n1062), .A1(n1395), .A2(n1074), .B0(n1046), .Y(n1394) );
  NOR2X1 U2319 ( .A(n1889), .B(\iexec_stage/BUS476[27] ), .Y(n1046) );
  NAND2X1 U2320 ( .A(n1396), .B(n1397), .Y(\iexec_stage/BUS476[27] ) );
  AOI222XL U2321 ( .A0(cop_addr_o[27]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[27]), .C0(BUS7101[27]), .C1(n1377), .Y(n1397) );
  AOI222XL U2322 ( .A0(\iexec_stage/BUS2332[27] ), .A1(n1378), .B0(BUS7231[27]), .B1(n1379), .C0(n1380), .C1(n45), .Y(n1396) );
  CLKINVX1 U2323 ( .A(n549), .Y(n1889) );
  OAI221X1 U2324 ( .A0(n1381), .A1(n1398), .B0(n1383), .B1(n1399), .C0(n1400), 
        .Y(n549) );
  AOI22X1 U2325 ( .A0(cop_addr_o[27]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[27]), .Y(n1400) );
  CLKINVX1 U2326 ( .A(BUS7231[27]), .Y(n1398) );
  NAND2X1 U2327 ( .A(n1892), .B(\iexec_stage/BUS476[25] ), .Y(n1074) );
  CLKINVX1 U2328 ( .A(n551), .Y(n1892) );
  OAI211X1 U2329 ( .A0(n1111), .A1(n1401), .B0(n1075), .C0(n1096), .Y(n1395)
         );
  NAND2X1 U2330 ( .A(n552), .B(n580), .Y(n1096) );
  CLKINVX1 U2331 ( .A(\iexec_stage/BUS476[24] ), .Y(n580) );
  NAND2X1 U2332 ( .A(n551), .B(n579), .Y(n1075) );
  CLKINVX1 U2333 ( .A(\iexec_stage/BUS476[25] ), .Y(n579) );
  NAND2X1 U2334 ( .A(n1402), .B(n1403), .Y(\iexec_stage/BUS476[25] ) );
  AOI222XL U2335 ( .A0(cop_addr_o[25]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[25]), .C0(BUS7101[25]), .C1(n1377), .Y(n1403) );
  AOI222XL U2336 ( .A0(\iexec_stage/BUS2332[25] ), .A1(n1378), .B0(BUS7231[25]), .B1(n1379), .C0(n1380), .C1(n46), .Y(n1402) );
  OAI221X1 U2337 ( .A0(n1381), .A1(n1404), .B0(n1383), .B1(n1405), .C0(n1406), 
        .Y(n551) );
  AOI22X1 U2338 ( .A0(cop_addr_o[25]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[25]), .Y(n1406) );
  CLKINVX1 U2339 ( .A(BUS7231[25]), .Y(n1404) );
  OAI31X1 U2340 ( .A0(n1133), .A1(n1407), .A2(n1110), .B0(n1095), .Y(n1401) );
  NAND2X1 U2341 ( .A(n1893), .B(\iexec_stage/BUS476[24] ), .Y(n1095) );
  NAND2X1 U2342 ( .A(n1408), .B(n1409), .Y(\iexec_stage/BUS476[24] ) );
  AOI222XL U2343 ( .A0(cop_addr_o[24]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[24]), .C0(BUS7101[24]), .C1(n1377), .Y(n1409) );
  AOI222XL U2344 ( .A0(\iexec_stage/BUS2332[24] ), .A1(n1378), .B0(BUS7231[24]), .B1(n1379), .C0(n1380), .C1(n47), .Y(n1408) );
  CLKINVX1 U2345 ( .A(n552), .Y(n1893) );
  OAI221X1 U2346 ( .A0(n1381), .A1(n1410), .B0(n1383), .B1(n1411), .C0(n1412), 
        .Y(n552) );
  CLKINVX1 U2347 ( .A(BUS7231[24]), .Y(n1410) );
  NOR2X1 U2348 ( .A(n1895), .B(\iexec_stage/BUS476[23] ), .Y(n1110) );
  CLKINVX1 U2349 ( .A(n553), .Y(n1895) );
  AOI211X1 U2350 ( .A0(n1413), .A1(n1163), .B0(n1146), .C0(n1132), .Y(n1407)
         );
  NOR2X1 U2351 ( .A(n554), .B(n582), .Y(n1132) );
  CLKINVX1 U2352 ( .A(\iexec_stage/BUS476[22] ), .Y(n582) );
  NOR2X1 U2353 ( .A(n555), .B(n583), .Y(n1146) );
  CLKINVX1 U2354 ( .A(\iexec_stage/BUS476[21] ), .Y(n583) );
  NAND2X1 U2355 ( .A(n556), .B(n584), .Y(n1163) );
  CLKINVX1 U2356 ( .A(\iexec_stage/BUS476[20] ), .Y(n584) );
  AOI31X1 U2357 ( .A0(n1162), .A1(n1414), .A2(n1189), .B0(n1145), .Y(n1413) );
  NOR2X1 U2358 ( .A(n1897), .B(\iexec_stage/BUS476[21] ), .Y(n1145) );
  NAND2X1 U2359 ( .A(n1415), .B(n1416), .Y(\iexec_stage/BUS476[21] ) );
  AOI222XL U2360 ( .A0(cop_addr_o[21]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[21]), .C0(BUS7101[21]), .C1(n1377), .Y(n1416) );
  AOI222XL U2361 ( .A0(\iexec_stage/BUS2332[21] ), .A1(n1378), .B0(BUS7231[21]), .B1(n1379), .C0(n1380), .C1(n48), .Y(n1415) );
  CLKINVX1 U2362 ( .A(n555), .Y(n1897) );
  OAI221X1 U2363 ( .A0(n1381), .A1(n1417), .B0(n1383), .B1(n1418), .C0(n1419), 
        .Y(n555) );
  CLKINVX1 U2364 ( .A(BUS7231[21]), .Y(n1417) );
  NAND2X1 U2365 ( .A(n1899), .B(\iexec_stage/BUS476[19] ), .Y(n1189) );
  CLKINVX1 U2366 ( .A(n557), .Y(n1899) );
  OAI211X1 U2367 ( .A0(n1224), .A1(n1420), .B0(n1188), .C0(n1206), .Y(n1414)
         );
  NAND2X1 U2368 ( .A(n558), .B(n587), .Y(n1206) );
  CLKINVX1 U2369 ( .A(\iexec_stage/BUS476[18] ), .Y(n587) );
  NAND2X1 U2370 ( .A(n557), .B(n586), .Y(n1188) );
  CLKINVX1 U2371 ( .A(\iexec_stage/BUS476[19] ), .Y(n586) );
  NAND2X1 U2372 ( .A(n1421), .B(n1422), .Y(\iexec_stage/BUS476[19] ) );
  AOI222XL U2373 ( .A0(cop_addr_o[19]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[19]), .C0(BUS7101[19]), .C1(n1377), .Y(n1422) );
  AOI222XL U2374 ( .A0(\iexec_stage/BUS2332[19] ), .A1(n1378), .B0(BUS7231[19]), .B1(n1379), .C0(n1380), .C1(n49), .Y(n1421) );
  OAI221X1 U2375 ( .A0(n1381), .A1(n1423), .B0(n1383), .B1(n1424), .C0(n1425), 
        .Y(n557) );
  CLKINVX1 U2376 ( .A(BUS7231[19]), .Y(n1423) );
  OAI31X1 U2377 ( .A0(n1242), .A1(n1426), .A2(n1223), .B0(n1205), .Y(n1420) );
  NAND2X1 U2378 ( .A(n1901), .B(\iexec_stage/BUS476[18] ), .Y(n1205) );
  NAND2X1 U2379 ( .A(n1427), .B(n1428), .Y(\iexec_stage/BUS476[18] ) );
  AOI222XL U2380 ( .A0(cop_addr_o[18]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[18]), .C0(BUS7101[18]), .C1(n1377), .Y(n1428) );
  AOI222XL U2381 ( .A0(\iexec_stage/BUS2332[18] ), .A1(n1378), .B0(BUS7231[18]), .B1(n1379), .C0(n1380), .C1(n50), .Y(n1427) );
  CLKINVX1 U2382 ( .A(n558), .Y(n1901) );
  OAI221X1 U2383 ( .A0(n1381), .A1(n1429), .B0(n1383), .B1(n1430), .C0(n1431), 
        .Y(n558) );
  CLKINVX1 U2384 ( .A(BUS7231[18]), .Y(n1429) );
  NOR2X1 U2385 ( .A(n1903), .B(\iexec_stage/BUS476[17] ), .Y(n1223) );
  CLKINVX1 U2386 ( .A(n559), .Y(n1903) );
  AOI211X1 U2387 ( .A0(n1432), .A1(n1282), .B0(n1260), .C0(n1241), .Y(n1426)
         );
  NOR2X1 U2388 ( .A(n567), .B(n589), .Y(n1241) );
  CLKINVX1 U2389 ( .A(\iexec_stage/BUS476[16] ), .Y(n589) );
  NOR2X1 U2390 ( .A(n590), .B(\iexec_stage/BUS468[15] ), .Y(n1260) );
  CLKINVX1 U2391 ( .A(\iexec_stage/BUS476[15] ), .Y(n590) );
  NAND2X1 U2392 ( .A(n560), .B(n591), .Y(n1282) );
  CLKINVX1 U2393 ( .A(\iexec_stage/BUS476[14] ), .Y(n591) );
  AOI31X1 U2394 ( .A0(n1283), .A1(n1433), .A2(n1301), .B0(n1261), .Y(n1432) );
  NOR2X1 U2395 ( .A(n1909), .B(\iexec_stage/BUS476[15] ), .Y(n1261) );
  NAND2X1 U2396 ( .A(n1434), .B(n1435), .Y(\iexec_stage/BUS476[15] ) );
  AOI222XL U2397 ( .A0(cop_addr_o[15]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[15]), .C0(BUS7101[15]), .C1(n1377), .Y(n1435) );
  AOI222XL U2398 ( .A0(\iexec_stage/BUS2332[15] ), .A1(n1378), .B0(BUS7231[15]), .B1(n1379), .C0(n1380), .C1(n51), .Y(n1434) );
  CLKINVX1 U2399 ( .A(\iexec_stage/BUS468[15] ), .Y(n1909) );
  OAI221X1 U2400 ( .A0(n1381), .A1(n1436), .B0(n1383), .B1(n1437), .C0(n1438), 
        .Y(\iexec_stage/BUS468[15] ) );
  CLKINVX1 U2401 ( .A(BUS7231[15]), .Y(n1436) );
  NAND2X1 U2402 ( .A(n1912), .B(\iexec_stage/BUS476[13] ), .Y(n1301) );
  CLKINVX1 U2403 ( .A(n561), .Y(n1912) );
  OAI211X1 U2404 ( .A0(n1335), .A1(n1439), .B0(n1302), .C0(n1319), .Y(n1433)
         );
  NAND2X1 U2405 ( .A(n562), .B(n593), .Y(n1319) );
  CLKINVX1 U2406 ( .A(\iexec_stage/BUS476[12] ), .Y(n593) );
  NAND2X1 U2407 ( .A(n561), .B(n592), .Y(n1302) );
  CLKINVX1 U2408 ( .A(\iexec_stage/BUS476[13] ), .Y(n592) );
  NAND2X1 U2409 ( .A(n1440), .B(n1441), .Y(\iexec_stage/BUS476[13] ) );
  AOI222XL U2410 ( .A0(cop_addr_o[13]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[13]), .C0(BUS7101[13]), .C1(n1377), .Y(n1441) );
  AOI222XL U2411 ( .A0(\iexec_stage/BUS2332[13] ), .A1(n1378), .B0(BUS7231[13]), .B1(n1379), .C0(n1380), .C1(n52), .Y(n1440) );
  OAI221X1 U2412 ( .A0(n1381), .A1(n1442), .B0(n1383), .B1(n1443), .C0(n1444), 
        .Y(n561) );
  CLKINVX1 U2413 ( .A(BUS7231[13]), .Y(n1442) );
  OAI31X1 U2414 ( .A0(n1352), .A1(n1445), .A2(n1336), .B0(n1320), .Y(n1439) );
  NAND2X1 U2415 ( .A(n1913), .B(\iexec_stage/BUS476[12] ), .Y(n1320) );
  NAND2X1 U2416 ( .A(n1446), .B(n1447), .Y(\iexec_stage/BUS476[12] ) );
  AOI222XL U2417 ( .A0(cop_addr_o[12]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[12]), .C0(BUS7101[12]), .C1(n1377), .Y(n1447) );
  AOI222XL U2418 ( .A0(\iexec_stage/BUS2332[12] ), .A1(n1378), .B0(BUS7231[12]), .B1(n1379), .C0(n1380), .C1(n53), .Y(n1446) );
  CLKINVX1 U2419 ( .A(n562), .Y(n1913) );
  OAI221X1 U2420 ( .A0(n1381), .A1(n1448), .B0(n1383), .B1(n1449), .C0(n1450), 
        .Y(n562) );
  CLKINVX1 U2421 ( .A(BUS7231[12]), .Y(n1448) );
  NOR2X1 U2422 ( .A(n1915), .B(\iexec_stage/BUS476[11] ), .Y(n1336) );
  CLKINVX1 U2423 ( .A(n563), .Y(n1915) );
  AOI211X1 U2424 ( .A0(n1451), .A1(n893), .B0(n1351), .C0(n866), .Y(n1445) );
  NOR2X1 U2425 ( .A(n568), .B(\iexec_stage/BUS468[9] ), .Y(n866) );
  CLKINVX1 U2426 ( .A(\iexec_stage/BUS476[9] ), .Y(n568) );
  NOR2X1 U2427 ( .A(n564), .B(n595), .Y(n1351) );
  CLKINVX1 U2428 ( .A(\iexec_stage/BUS476[10] ), .Y(n595) );
  NAND2X1 U2429 ( .A(n539), .B(n569), .Y(n893) );
  CLKINVX1 U2430 ( .A(\iexec_stage/BUS476[8] ), .Y(n569) );
  AOI31X1 U2431 ( .A0(n894), .A1(n1452), .A2(n914), .B0(n867), .Y(n1451) );
  NOR2X1 U2432 ( .A(n1917), .B(\iexec_stage/BUS476[9] ), .Y(n867) );
  NAND2X1 U2433 ( .A(n1453), .B(n1454), .Y(\iexec_stage/BUS476[9] ) );
  AOI222XL U2434 ( .A0(cop_addr_o[9]), .A1(n1375), .B0(n1376), .B1(BUS15471[9]), .C0(BUS7101[9]), .C1(n1377), .Y(n1454) );
  AOI222XL U2435 ( .A0(\iexec_stage/BUS2332[9] ), .A1(n1378), .B0(BUS7231[9]), 
        .B1(n1379), .C0(n1380), .C1(n54), .Y(n1453) );
  CLKINVX1 U2436 ( .A(\iexec_stage/BUS468[9] ), .Y(n1917) );
  OAI221X1 U2437 ( .A0(n1381), .A1(n1455), .B0(n1383), .B1(n1456), .C0(n1457), 
        .Y(\iexec_stage/BUS468[9] ) );
  AOI22X1 U2438 ( .A0(cop_addr_o[9]), .A1(n1386), .B0(n1387), .B1(BUS15471[9]), 
        .Y(n1457) );
  CLKINVX1 U2439 ( .A(BUS7231[9]), .Y(n1455) );
  NAND2X1 U2440 ( .A(n1919), .B(\iexec_stage/BUS476[7] ), .Y(n914) );
  CLKINVX1 U2441 ( .A(n540), .Y(n1919) );
  OAI211X1 U2442 ( .A0(n941), .A1(n1458), .B0(n915), .C0(n928), .Y(n1452) );
  NAND2X1 U2443 ( .A(n541), .B(n571), .Y(n928) );
  CLKINVX1 U2444 ( .A(\iexec_stage/BUS476[6] ), .Y(n571) );
  NAND2X1 U2445 ( .A(n540), .B(n570), .Y(n915) );
  CLKINVX1 U2446 ( .A(\iexec_stage/BUS476[7] ), .Y(n570) );
  NAND2X1 U2447 ( .A(n1459), .B(n1460), .Y(\iexec_stage/BUS476[7] ) );
  AOI222XL U2448 ( .A0(cop_addr_o[7]), .A1(n1375), .B0(n1376), .B1(BUS15471[7]), .C0(BUS7101[7]), .C1(n1377), .Y(n1460) );
  AOI222XL U2449 ( .A0(\iexec_stage/BUS2332[7] ), .A1(n1378), .B0(BUS7231[7]), 
        .B1(n1379), .C0(n1380), .C1(n55), .Y(n1459) );
  OAI221X1 U2450 ( .A0(n1381), .A1(n1461), .B0(n1383), .B1(n720), .C0(n1462), 
        .Y(n540) );
  CLKINVX1 U2451 ( .A(BUS7117[7]), .Y(n720) );
  CLKINVX1 U2452 ( .A(BUS7231[7]), .Y(n1461) );
  OAI31X1 U2453 ( .A0(n954), .A1(n1463), .A2(n942), .B0(n929), .Y(n1458) );
  NAND2X1 U2454 ( .A(n1920), .B(\iexec_stage/BUS476[6] ), .Y(n929) );
  NAND2X1 U2455 ( .A(n1464), .B(n1465), .Y(\iexec_stage/BUS476[6] ) );
  AOI222XL U2456 ( .A0(cop_addr_o[6]), .A1(n1375), .B0(n1376), .B1(BUS15471[6]), .C0(BUS7101[6]), .C1(n1377), .Y(n1465) );
  AOI222XL U2457 ( .A0(\iexec_stage/BUS2332[6] ), .A1(n1378), .B0(BUS7231[6]), 
        .B1(n1379), .C0(n1380), .C1(n56), .Y(n1464) );
  CLKINVX1 U2458 ( .A(n541), .Y(n1920) );
  OAI221X1 U2459 ( .A0(n1381), .A1(n1466), .B0(n1383), .B1(n723), .C0(n1467), 
        .Y(n541) );
  AOI22X1 U2460 ( .A0(cop_addr_o[6]), .A1(n1386), .B0(n1387), .B1(BUS15471[6]), 
        .Y(n1467) );
  CLKINVX1 U2461 ( .A(BUS7117[6]), .Y(n723) );
  CLKINVX1 U2462 ( .A(BUS7231[6]), .Y(n1466) );
  NOR2X1 U2463 ( .A(n1921), .B(\iexec_stage/BUS476[5] ), .Y(n942) );
  CLKINVX1 U2464 ( .A(n542), .Y(n1921) );
  AOI211X1 U2465 ( .A0(n1468), .A1(n1001), .B0(n964), .C0(n955), .Y(n1463) );
  NOR2X1 U2466 ( .A(n543), .B(n1923), .Y(n955) );
  NOR2X1 U2467 ( .A(n544), .B(n574), .Y(n964) );
  NAND2X1 U2468 ( .A(n546), .B(n585), .Y(n1001) );
  AOI31X1 U2469 ( .A0(n1002), .A1(n1469), .A2(n1470), .B0(n965), .Y(n1468) );
  NOR2X1 U2470 ( .A(n1924), .B(\iexec_stage/BUS476[3] ), .Y(n965) );
  CLKINVX1 U2471 ( .A(n544), .Y(n1924) );
  OAI221X1 U2472 ( .A0(n1381), .A1(n1471), .B0(n1383), .B1(n732), .C0(n1472), 
        .Y(n544) );
  CLKINVX1 U2473 ( .A(BUS7117[3]), .Y(n732) );
  CLKINVX1 U2474 ( .A(BUS7231[3]), .Y(n1471) );
  CLKINVX1 U2475 ( .A(\iexec_stage/BUS468[1] ), .Y(n1926) );
  OAI221X1 U2476 ( .A0(n1381), .A1(n1473), .B0(n1383), .B1(n716), .C0(n1474), 
        .Y(\iexec_stage/BUS468[1] ) );
  AOI22X1 U2477 ( .A0(cop_addr_o[1]), .A1(n1386), .B0(n1387), .B1(BUS15471[1]), 
        .Y(n1474) );
  CLKINVX1 U2478 ( .A(BUS7117[1]), .Y(n716) );
  CLKINVX1 U2479 ( .A(BUS7231[1]), .Y(n1473) );
  CLKINVX1 U2480 ( .A(n546), .Y(n1925) );
  OAI221X1 U2481 ( .A0(n1381), .A1(n1475), .B0(n1383), .B1(n735), .C0(n1476), 
        .Y(n546) );
  CLKINVX1 U2482 ( .A(BUS7117[2]), .Y(n735) );
  CLKINVX1 U2483 ( .A(BUS7231[2]), .Y(n1475) );
  NOR2X1 U2484 ( .A(n1922), .B(\iexec_stage/BUS476[4] ), .Y(n954) );
  CLKINVX1 U2485 ( .A(n543), .Y(n1922) );
  OAI221X1 U2486 ( .A0(n1381), .A1(n1477), .B0(n1383), .B1(n729), .C0(n1478), 
        .Y(n543) );
  AOI22X1 U2487 ( .A0(cop_addr_o[4]), .A1(n1386), .B0(n1387), .B1(BUS15471[4]), 
        .Y(n1478) );
  CLKINVX1 U2488 ( .A(BUS7117[4]), .Y(n729) );
  CLKINVX1 U2489 ( .A(BUS7231[4]), .Y(n1477) );
  NOR2X1 U2490 ( .A(n542), .B(n572), .Y(n941) );
  CLKINVX1 U2491 ( .A(\iexec_stage/BUS476[5] ), .Y(n572) );
  NAND2X1 U2492 ( .A(n1479), .B(n1480), .Y(\iexec_stage/BUS476[5] ) );
  AOI222XL U2493 ( .A0(cop_addr_o[5]), .A1(n1375), .B0(n1376), .B1(BUS15471[5]), .C0(BUS7101[5]), .C1(n1377), .Y(n1480) );
  AOI222XL U2494 ( .A0(\iexec_stage/BUS2332[5] ), .A1(n1378), .B0(BUS7231[5]), 
        .B1(n1379), .C0(n1380), .C1(n57), .Y(n1479) );
  OAI221X1 U2495 ( .A0(n1381), .A1(n1481), .B0(n1383), .B1(n726), .C0(n1482), 
        .Y(n542) );
  AOI22X1 U2496 ( .A0(cop_addr_o[5]), .A1(n1386), .B0(n1387), .B1(BUS15471[5]), 
        .Y(n1482) );
  CLKINVX1 U2497 ( .A(BUS7117[5]), .Y(n726) );
  CLKINVX1 U2498 ( .A(BUS7231[5]), .Y(n1481) );
  NAND2X1 U2499 ( .A(n1918), .B(\iexec_stage/BUS476[8] ), .Y(n894) );
  NAND2X1 U2500 ( .A(n1483), .B(n1484), .Y(\iexec_stage/BUS476[8] ) );
  AOI222XL U2501 ( .A0(cop_addr_o[8]), .A1(n1375), .B0(n1376), .B1(BUS15471[8]), .C0(BUS7101[8]), .C1(n1377), .Y(n1484) );
  AOI222XL U2502 ( .A0(\iexec_stage/BUS2332[8] ), .A1(n1378), .B0(BUS7231[8]), 
        .B1(n1379), .C0(n1380), .C1(n58), .Y(n1483) );
  CLKINVX1 U2503 ( .A(n539), .Y(n1918) );
  OAI221X1 U2504 ( .A0(n1381), .A1(n1485), .B0(n1383), .B1(n1486), .C0(n1487), 
        .Y(n539) );
  CLKINVX1 U2505 ( .A(BUS7231[8]), .Y(n1485) );
  NOR2X1 U2506 ( .A(n1916), .B(\iexec_stage/BUS476[10] ), .Y(n1352) );
  NAND2X1 U2507 ( .A(n1488), .B(n1489), .Y(\iexec_stage/BUS476[10] ) );
  AOI222XL U2508 ( .A0(cop_addr_o[10]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[10]), .C0(BUS7101[10]), .C1(n1377), .Y(n1489) );
  AOI222XL U2509 ( .A0(\iexec_stage/BUS2332[10] ), .A1(n1378), .B0(BUS7231[10]), .B1(n1379), .C0(n1380), .C1(n59), .Y(n1488) );
  CLKINVX1 U2510 ( .A(n564), .Y(n1916) );
  OAI221X1 U2511 ( .A0(n1381), .A1(n1490), .B0(n1383), .B1(n1491), .C0(n1492), 
        .Y(n564) );
  CLKINVX1 U2512 ( .A(BUS7231[10]), .Y(n1490) );
  NOR2X1 U2513 ( .A(n563), .B(n594), .Y(n1335) );
  CLKINVX1 U2514 ( .A(\iexec_stage/BUS476[11] ), .Y(n594) );
  NAND2X1 U2515 ( .A(n1493), .B(n1494), .Y(\iexec_stage/BUS476[11] ) );
  AOI222XL U2516 ( .A0(cop_addr_o[11]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[11]), .C0(BUS7101[11]), .C1(n1377), .Y(n1494) );
  AOI222XL U2517 ( .A0(\iexec_stage/BUS2332[11] ), .A1(n1378), .B0(BUS7231[11]), .B1(n1379), .C0(n1380), .C1(n60), .Y(n1493) );
  OAI221X1 U2518 ( .A0(n1381), .A1(n1495), .B0(n1383), .B1(n1496), .C0(n1497), 
        .Y(n563) );
  CLKINVX1 U2519 ( .A(BUS7231[11]), .Y(n1495) );
  NAND2X1 U2520 ( .A(n1911), .B(\iexec_stage/BUS476[14] ), .Y(n1283) );
  NAND2X1 U2521 ( .A(n1498), .B(n1499), .Y(\iexec_stage/BUS476[14] ) );
  AOI222XL U2522 ( .A0(cop_addr_o[14]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[14]), .C0(BUS7101[14]), .C1(n1377), .Y(n1499) );
  AOI222XL U2523 ( .A0(\iexec_stage/BUS2332[14] ), .A1(n1378), .B0(BUS7231[14]), .B1(n1379), .C0(n1380), .C1(n61), .Y(n1498) );
  CLKINVX1 U2524 ( .A(n560), .Y(n1911) );
  OAI221X1 U2525 ( .A0(n1381), .A1(n1500), .B0(n1383), .B1(n1501), .C0(n1502), 
        .Y(n560) );
  CLKINVX1 U2526 ( .A(BUS7231[14]), .Y(n1500) );
  NOR2X1 U2527 ( .A(n1906), .B(\iexec_stage/BUS476[16] ), .Y(n1242) );
  NAND2X1 U2528 ( .A(n1503), .B(n1504), .Y(\iexec_stage/BUS476[16] ) );
  AOI222XL U2529 ( .A0(cop_addr_o[16]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[16]), .C0(BUS7101[16]), .C1(n1377), .Y(n1504) );
  AOI222XL U2530 ( .A0(\iexec_stage/BUS2332[16] ), .A1(n1378), .B0(BUS7231[16]), .B1(n1379), .C0(n1380), .C1(n62), .Y(n1503) );
  CLKINVX1 U2531 ( .A(n567), .Y(n1906) );
  OAI221X1 U2532 ( .A0(n1381), .A1(n1505), .B0(n1383), .B1(n1506), .C0(n1507), 
        .Y(n567) );
  CLKINVX1 U2533 ( .A(BUS7231[16]), .Y(n1505) );
  NOR2X1 U2534 ( .A(n559), .B(n588), .Y(n1224) );
  CLKINVX1 U2535 ( .A(\iexec_stage/BUS476[17] ), .Y(n588) );
  NAND2X1 U2536 ( .A(n1508), .B(n1509), .Y(\iexec_stage/BUS476[17] ) );
  AOI222XL U2537 ( .A0(cop_addr_o[17]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[17]), .C0(BUS7101[17]), .C1(n1377), .Y(n1509) );
  AOI222XL U2538 ( .A0(\iexec_stage/BUS2332[17] ), .A1(n1378), .B0(BUS7231[17]), .B1(n1379), .C0(n1380), .C1(n63), .Y(n1508) );
  OAI221X1 U2539 ( .A0(n1381), .A1(n1510), .B0(n1383), .B1(n1511), .C0(n1512), 
        .Y(n559) );
  CLKINVX1 U2540 ( .A(BUS7231[17]), .Y(n1510) );
  NAND2X1 U2541 ( .A(n1898), .B(\iexec_stage/BUS476[20] ), .Y(n1162) );
  NAND2X1 U2542 ( .A(n1513), .B(n1514), .Y(\iexec_stage/BUS476[20] ) );
  AOI222XL U2543 ( .A0(cop_addr_o[20]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[20]), .C0(BUS7101[20]), .C1(n1377), .Y(n1514) );
  AOI222XL U2544 ( .A0(\iexec_stage/BUS2332[20] ), .A1(n1378), .B0(BUS7231[20]), .B1(n1379), .C0(n1380), .C1(n64), .Y(n1513) );
  CLKINVX1 U2545 ( .A(n556), .Y(n1898) );
  OAI221X1 U2546 ( .A0(n1381), .A1(n1515), .B0(n1383), .B1(n1516), .C0(n1517), 
        .Y(n556) );
  CLKINVX1 U2547 ( .A(BUS7231[20]), .Y(n1515) );
  NOR2X1 U2548 ( .A(n1896), .B(\iexec_stage/BUS476[22] ), .Y(n1133) );
  NAND2X1 U2549 ( .A(n1518), .B(n1519), .Y(\iexec_stage/BUS476[22] ) );
  AOI222XL U2550 ( .A0(cop_addr_o[22]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[22]), .C0(BUS7101[22]), .C1(n1377), .Y(n1519) );
  AOI222XL U2551 ( .A0(\iexec_stage/BUS2332[22] ), .A1(n1378), .B0(BUS7231[22]), .B1(n1379), .C0(n1380), .C1(n65), .Y(n1518) );
  CLKINVX1 U2552 ( .A(n554), .Y(n1896) );
  OAI221X1 U2553 ( .A0(n1381), .A1(n1520), .B0(n1383), .B1(n1521), .C0(n1522), 
        .Y(n554) );
  CLKINVX1 U2554 ( .A(BUS7231[22]), .Y(n1520) );
  NOR2X1 U2555 ( .A(n553), .B(n581), .Y(n1111) );
  CLKINVX1 U2556 ( .A(\iexec_stage/BUS476[23] ), .Y(n581) );
  NAND2X1 U2557 ( .A(n1523), .B(n1524), .Y(\iexec_stage/BUS476[23] ) );
  AOI222XL U2558 ( .A0(cop_addr_o[23]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[23]), .C0(BUS7101[23]), .C1(n1377), .Y(n1524) );
  AOI222XL U2559 ( .A0(\iexec_stage/BUS2332[23] ), .A1(n1378), .B0(BUS7231[23]), .B1(n1379), .C0(n1380), .C1(n66), .Y(n1523) );
  OAI221X1 U2560 ( .A0(n1381), .A1(n1525), .B0(n1383), .B1(n1526), .C0(n1527), 
        .Y(n553) );
  AOI22X1 U2561 ( .A0(cop_addr_o[23]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[23]), .Y(n1527) );
  CLKINVX1 U2562 ( .A(BUS7231[23]), .Y(n1525) );
  NAND2X1 U2563 ( .A(n1891), .B(\iexec_stage/BUS476[26] ), .Y(n1062) );
  NAND2X1 U2564 ( .A(n1528), .B(n1529), .Y(\iexec_stage/BUS476[26] ) );
  AOI222XL U2565 ( .A0(cop_addr_o[26]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[26]), .C0(BUS7101[26]), .C1(n1377), .Y(n1529) );
  AOI222XL U2566 ( .A0(\iexec_stage/BUS2332[26] ), .A1(n1378), .B0(BUS7231[26]), .B1(n1379), .C0(n1380), .C1(n67), .Y(n1528) );
  CLKINVX1 U2567 ( .A(n550), .Y(n1891) );
  OAI221X1 U2568 ( .A0(n1381), .A1(n1530), .B0(n1383), .B1(n1531), .C0(n1532), 
        .Y(n550) );
  AOI22X1 U2569 ( .A0(cop_addr_o[26]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[26]), .Y(n1532) );
  CLKINVX1 U2570 ( .A(BUS7231[26]), .Y(n1530) );
  NOR2X1 U2571 ( .A(n1886), .B(\iexec_stage/BUS476[28] ), .Y(n1035) );
  NAND2X1 U2572 ( .A(n1533), .B(n1534), .Y(\iexec_stage/BUS476[28] ) );
  AOI222XL U2573 ( .A0(cop_addr_o[28]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[28]), .C0(BUS7101[28]), .C1(n1377), .Y(n1534) );
  AOI222XL U2574 ( .A0(\iexec_stage/BUS2332[28] ), .A1(n1378), .B0(BUS7231[28]), .B1(n1379), .C0(n1380), .C1(n73), .Y(n1533) );
  CLKINVX1 U2575 ( .A(n548), .Y(n1886) );
  OAI221X1 U2576 ( .A0(n1381), .A1(n1535), .B0(n1383), .B1(n1536), .C0(n1537), 
        .Y(n548) );
  AOI22X1 U2577 ( .A0(cop_addr_o[28]), .A1(n1386), .B0(n1387), .B1(
        BUS15471[28]), .Y(n1537) );
  CLKINVX1 U2578 ( .A(BUS7231[28]), .Y(n1535) );
  CLKINVX1 U2579 ( .A(\iexec_stage/BUS468[31] ), .Y(n1881) );
  OAI221X1 U2580 ( .A0(n1381), .A1(n1538), .B0(n1383), .B1(n1539), .C0(n1540), 
        .Y(\iexec_stage/BUS468[31] ) );
  CLKINVX1 U2581 ( .A(BUS7231[31]), .Y(n1538) );
  NAND2X1 U2582 ( .A(n1541), .B(n1542), .Y(\iexec_stage/BUS476[31] ) );
  AOI222XL U2583 ( .A0(cop_addr_o[31]), .A1(n1375), .B0(n1376), .B1(
        BUS15471[31]), .C0(BUS7101[31]), .C1(n1377), .Y(n1542) );
  AOI222XL U2584 ( .A0(\iexec_stage/BUS2332[31] ), .A1(n1378), .B0(BUS7231[31]), .B1(n1379), .C0(n1380), .C1(n74), .Y(n1541) );
  CLKINVX1 U2585 ( .A(n967), .Y(n889) );
  AOI2BB1X1 U2586 ( .A0N(n951), .A1N(n980), .B0(n857), .Y(n967) );
  CLKINVX1 U2587 ( .A(n982), .Y(n857) );
  MXI2X1 U2588 ( .A(n1543), .B(n862), .S0(n286), .Y(n982) );
  NOR2X1 U2589 ( .A(n287), .B(n1544), .Y(n1543) );
  NAND2X1 U2590 ( .A(n1358), .B(n1360), .Y(n980) );
  NOR2X1 U2591 ( .A(\iexec_stage/BUS476[1] ), .B(\iexec_stage/BUS476[3] ), .Y(
        n1360) );
  AOI222XL U2592 ( .A0(cop_addr_o[3]), .A1(n1375), .B0(n1376), .B1(BUS15471[3]), .C0(BUS7101[3]), .C1(n1377), .Y(n1546) );
  AOI222XL U2593 ( .A0(\iexec_stage/BUS2332[3] ), .A1(n1378), .B0(BUS7231[3]), 
        .B1(n1379), .C0(n1380), .C1(n68), .Y(n1545) );
  AOI222XL U2594 ( .A0(cop_addr_o[1]), .A1(n1375), .B0(n1376), .B1(BUS15471[1]), .C0(BUS7101[1]), .C1(n1377), .Y(n1548) );
  AOI222XL U2595 ( .A0(\iexec_stage/BUS2332[1] ), .A1(n1378), .B0(BUS7231[1]), 
        .B1(n1379), .C0(n1380), .C1(n75), .Y(n1547) );
  AND2X1 U2596 ( .A(n1362), .B(n585), .Y(n1358) );
  AOI222XL U2597 ( .A0(cop_addr_o[2]), .A1(n1375), .B0(n1376), .B1(BUS15471[2]), .C0(BUS7101[2]), .C1(n1377), .Y(n1550) );
  AOI222XL U2598 ( .A0(\iexec_stage/BUS2332[2] ), .A1(n1378), .B0(BUS7231[2]), 
        .B1(n1379), .C0(n1380), .C1(n69), .Y(n1549) );
  NOR2X1 U2599 ( .A(\iexec_stage/BUS476[0] ), .B(\iexec_stage/BUS476[4] ), .Y(
        n1362) );
  AOI222XL U2600 ( .A0(cop_addr_o[4]), .A1(n1375), .B0(n1376), .B1(BUS15471[4]), .C0(BUS7101[4]), .C1(n1377), .Y(n1552) );
  AOI222XL U2601 ( .A0(\iexec_stage/BUS2332[4] ), .A1(n1378), .B0(BUS7231[4]), 
        .B1(n1379), .C0(n1380), .C1(n70), .Y(n1551) );
  NAND2X1 U2602 ( .A(n1031), .B(n1024), .Y(n951) );
  CLKINVX1 U2603 ( .A(n1043), .Y(n1024) );
  NAND2X1 U2604 ( .A(n290), .B(n289), .Y(n1043) );
  NOR3BX1 U2605 ( .AN(n288), .B(n40), .C(n287), .Y(n1031) );
  AOI221XL U2606 ( .A0(\iexec_stage/MIPS_alu/mips_alu/N370 ), .A1(n1938), .B0(
        \iexec_stage/MIPS_alu/mips_alu/N112 ), .B1(n855), .C0(n1553), .Y(n1363) );
  MXI2X1 U2607 ( .A(n1554), .B(n1555), .S0(n597), .Y(n1553) );
  AOI222XL U2608 ( .A0(n1375), .A1(cop_addr_o[0]), .B0(n1376), .B1(BUS15471[0]), .C0(BUS7101[0]), .C1(n1377), .Y(n1557) );
  AND3X2 U2609 ( .A(n1558), .B(n1559), .C(n1560), .Y(n1377) );
  AND3X2 U2610 ( .A(n1561), .B(n1559), .C(n1560), .Y(n1376) );
  CLKINVX1 U2611 ( .A(n1558), .Y(n1561) );
  NAND4X1 U2612 ( .A(n1562), .B(n1563), .C(n1564), .D(n1565), .Y(n1558) );
  NOR3X1 U2613 ( .A(n1566), .B(n1567), .C(n1568), .Y(n1565) );
  XOR2X1 U2614 ( .A(\iforward/BUS82[2] ), .B(BUS18211[2]), .Y(n1568) );
  XOR2X1 U2615 ( .A(\iforward/BUS82[4] ), .B(BUS18211[4]), .Y(n1567) );
  XOR2X1 U2616 ( .A(\iforward/BUS82[3] ), .B(BUS18211[3]), .Y(n1566) );
  XOR2X1 U2617 ( .A(\iforward/BUS82[0] ), .B(n1569), .Y(n1564) );
  XOR2X1 U2618 ( .A(\iforward/BUS82[1] ), .B(n1570), .Y(n1562) );
  NOR2BX1 U2619 ( .AN(n1560), .B(n1559), .Y(n1375) );
  NAND4X1 U2620 ( .A(n1571), .B(n1572), .C(n1573), .D(n1574), .Y(n1559) );
  NOR3X1 U2621 ( .A(n1575), .B(n1576), .C(n1577), .Y(n1574) );
  XOR2X1 U2622 ( .A(\iforward/BUS82[2] ), .B(BUS1724[2]), .Y(n1577) );
  XOR2X1 U2623 ( .A(\iforward/BUS82[4] ), .B(BUS1724[4]), .Y(n1576) );
  XOR2X1 U2624 ( .A(\iforward/BUS82[3] ), .B(BUS1724[3]), .Y(n1575) );
  XOR2X1 U2625 ( .A(\iforward/BUS82[0] ), .B(n1578), .Y(n1573) );
  XOR2X1 U2626 ( .A(\iforward/BUS82[1] ), .B(n1579), .Y(n1571) );
  AND2X1 U2627 ( .A(n291), .B(n77), .Y(n1560) );
  AOI222XL U2628 ( .A0(\iexec_stage/BUS2332[0] ), .A1(n1378), .B0(n1379), .B1(
        BUS7231[0]), .C0(n1380), .C1(n76), .Y(n1556) );
  AND2X1 U2629 ( .A(n292), .B(n291), .Y(n1380) );
  NOR2X1 U2630 ( .A(n291), .B(n292), .Y(n1379) );
  NOR2X1 U2631 ( .A(n77), .B(n291), .Y(n1378) );
  MXI2X1 U2632 ( .A(n868), .B(n978), .S0(n1927), .Y(n1555) );
  NOR3X1 U2633 ( .A(n1544), .B(n286), .C(n39), .Y(n978) );
  NOR2X1 U2634 ( .A(n979), .B(n1580), .Y(n1554) );
  MXI2X1 U2635 ( .A(n995), .B(n953), .S0(n1927), .Y(n1580) );
  CLKINVX1 U2636 ( .A(n565), .Y(n1927) );
  OAI221X1 U2637 ( .A0(n1381), .A1(n1581), .B0(n1383), .B1(n738), .C0(n1582), 
        .Y(n565) );
  AOI22X1 U2638 ( .A0(cop_addr_o[0]), .A1(n1386), .B0(n1387), .B1(BUS15471[0]), 
        .Y(n1582) );
  NOR3BX1 U2639 ( .AN(n281), .B(n280), .C(n714), .Y(n1387) );
  NOR3BX1 U2640 ( .AN(n281), .B(n711), .C(n280), .Y(n1386) );
  CLKINVX1 U2641 ( .A(BUS7117[0]), .Y(n738) );
  MXI2X1 U2642 ( .A(n1583), .B(n281), .S0(n280), .Y(n1383) );
  OAI2BB1X1 U2643 ( .A0N(n711), .A1N(n714), .B0(n281), .Y(n1583) );
  CLKINVX1 U2644 ( .A(BUS7231[0]), .Y(n1581) );
  NAND2BX1 U2645 ( .AN(n281), .B(n280), .Y(n1381) );
  CLKINVX1 U2646 ( .A(n868), .Y(n953) );
  NOR2X1 U2647 ( .A(n1366), .B(n1544), .Y(n868) );
  CLKINVX1 U2648 ( .A(n863), .Y(n979) );
  OAI2BB1X1 U2649 ( .A0N(n995), .A1N(n1584), .B0(n286), .Y(n863) );
  OR2X1 U2650 ( .A(n1544), .B(n287), .Y(n1584) );
  NAND3BX1 U2651 ( .AN(n288), .B(n289), .C(n36), .Y(n1544) );
  CLKINVX1 U2652 ( .A(n862), .Y(n995) );
  NOR2X1 U2653 ( .A(n1368), .B(n287), .Y(n862) );
  NOR3X1 U2654 ( .A(n36), .B(n289), .C(n1369), .Y(n855) );
  CLKINVX1 U2655 ( .A(n1078), .Y(n1369) );
  NOR2X1 U2656 ( .A(n1366), .B(n288), .Y(n1078) );
  NAND2X1 U2657 ( .A(n287), .B(n286), .Y(n1366) );
  NOR3X1 U2658 ( .A(n1368), .B(n286), .C(n39), .Y(n1938) );
  NAND3X1 U2659 ( .A(n288), .B(n36), .C(n289), .Y(n1368) );
  OAI222X1 U2660 ( .A0(n711), .A1(n1585), .B0(n1586), .B1(n714), .C0(n715), 
        .C1(n1456), .Y(BUS9884[9]) );
  CLKINVX1 U2661 ( .A(BUS7117[9]), .Y(n1456) );
  OAI222X1 U2662 ( .A0(n711), .A1(n1587), .B0(n1588), .B1(n714), .C0(n715), 
        .C1(n1486), .Y(BUS9884[8]) );
  CLKINVX1 U2663 ( .A(BUS7117[8]), .Y(n1486) );
  OAI222X1 U2664 ( .A0(n711), .A1(n1589), .B0(n1590), .B1(n714), .C0(n715), 
        .C1(n1539), .Y(BUS9884[31]) );
  CLKINVX1 U2665 ( .A(BUS7117[31]), .Y(n1539) );
  OAI222X1 U2666 ( .A0(n711), .A1(n1591), .B0(n1592), .B1(n714), .C0(n715), 
        .C1(n1384), .Y(BUS9884[30]) );
  CLKINVX1 U2667 ( .A(BUS7117[30]), .Y(n1384) );
  OAI222X1 U2668 ( .A0(n711), .A1(n1593), .B0(n1594), .B1(n714), .C0(n715), 
        .C1(n1392), .Y(BUS9884[29]) );
  CLKINVX1 U2669 ( .A(BUS7117[29]), .Y(n1392) );
  OAI222X1 U2670 ( .A0(n711), .A1(n1595), .B0(n1596), .B1(n714), .C0(n715), 
        .C1(n1536), .Y(BUS9884[28]) );
  CLKINVX1 U2671 ( .A(BUS7117[28]), .Y(n1536) );
  OAI222X1 U2672 ( .A0(n711), .A1(n1597), .B0(n1598), .B1(n714), .C0(n715), 
        .C1(n1399), .Y(BUS9884[27]) );
  CLKINVX1 U2673 ( .A(BUS7117[27]), .Y(n1399) );
  OAI222X1 U2674 ( .A0(n711), .A1(n1599), .B0(n1600), .B1(n714), .C0(n715), 
        .C1(n1531), .Y(BUS9884[26]) );
  CLKINVX1 U2675 ( .A(BUS7117[26]), .Y(n1531) );
  OAI222X1 U2676 ( .A0(n711), .A1(n1601), .B0(n1602), .B1(n714), .C0(n715), 
        .C1(n1405), .Y(BUS9884[25]) );
  CLKINVX1 U2677 ( .A(BUS7117[25]), .Y(n1405) );
  OAI222X1 U2678 ( .A0(n711), .A1(n1603), .B0(n1604), .B1(n714), .C0(n715), 
        .C1(n1411), .Y(BUS9884[24]) );
  CLKINVX1 U2679 ( .A(BUS7117[24]), .Y(n1411) );
  OAI222X1 U2680 ( .A0(n711), .A1(n1605), .B0(n1606), .B1(n714), .C0(n715), 
        .C1(n1526), .Y(BUS9884[23]) );
  CLKINVX1 U2681 ( .A(BUS7117[23]), .Y(n1526) );
  OAI222X1 U2682 ( .A0(n711), .A1(n1607), .B0(n1608), .B1(n714), .C0(n715), 
        .C1(n1521), .Y(BUS9884[22]) );
  CLKINVX1 U2683 ( .A(BUS7117[22]), .Y(n1521) );
  OAI222X1 U2684 ( .A0(n711), .A1(n1609), .B0(n1610), .B1(n714), .C0(n715), 
        .C1(n1418), .Y(BUS9884[21]) );
  CLKINVX1 U2685 ( .A(BUS7117[21]), .Y(n1418) );
  OAI222X1 U2686 ( .A0(n711), .A1(n1611), .B0(n1612), .B1(n714), .C0(n715), 
        .C1(n1516), .Y(BUS9884[20]) );
  CLKINVX1 U2687 ( .A(BUS7117[20]), .Y(n1516) );
  OAI222X1 U2688 ( .A0(n711), .A1(n1613), .B0(n1614), .B1(n714), .C0(n715), 
        .C1(n1424), .Y(BUS9884[19]) );
  CLKINVX1 U2689 ( .A(BUS7117[19]), .Y(n1424) );
  OAI222X1 U2690 ( .A0(n711), .A1(n1615), .B0(n1616), .B1(n714), .C0(n715), 
        .C1(n1430), .Y(BUS9884[18]) );
  CLKINVX1 U2691 ( .A(BUS7117[18]), .Y(n1430) );
  OAI222X1 U2692 ( .A0(n711), .A1(n1617), .B0(n1618), .B1(n714), .C0(n715), 
        .C1(n1511), .Y(BUS9884[17]) );
  CLKINVX1 U2693 ( .A(BUS7117[17]), .Y(n1511) );
  OAI222X1 U2694 ( .A0(n711), .A1(n1619), .B0(n1620), .B1(n714), .C0(n715), 
        .C1(n1506), .Y(BUS9884[16]) );
  CLKINVX1 U2695 ( .A(BUS7117[16]), .Y(n1506) );
  OAI222X1 U2696 ( .A0(n711), .A1(n1621), .B0(n1622), .B1(n714), .C0(n715), 
        .C1(n1437), .Y(BUS9884[15]) );
  CLKINVX1 U2697 ( .A(BUS7117[15]), .Y(n1437) );
  OAI222X1 U2698 ( .A0(n711), .A1(n1623), .B0(n1624), .B1(n714), .C0(n715), 
        .C1(n1501), .Y(BUS9884[14]) );
  CLKINVX1 U2699 ( .A(BUS7117[14]), .Y(n1501) );
  OAI222X1 U2700 ( .A0(n711), .A1(n1625), .B0(n1626), .B1(n714), .C0(n715), 
        .C1(n1443), .Y(BUS9884[13]) );
  CLKINVX1 U2701 ( .A(BUS7117[13]), .Y(n1443) );
  OAI222X1 U2702 ( .A0(n711), .A1(n1627), .B0(n1628), .B1(n714), .C0(n715), 
        .C1(n1449), .Y(BUS9884[12]) );
  CLKINVX1 U2703 ( .A(BUS7117[12]), .Y(n1449) );
  OAI222X1 U2704 ( .A0(n711), .A1(n1629), .B0(n1630), .B1(n714), .C0(n715), 
        .C1(n1496), .Y(BUS9884[11]) );
  CLKINVX1 U2705 ( .A(BUS7117[11]), .Y(n1496) );
  OAI222X1 U2706 ( .A0(n711), .A1(n1631), .B0(n1632), .B1(n714), .C0(n715), 
        .C1(n1491), .Y(BUS9884[10]) );
  CLKINVX1 U2707 ( .A(BUS7117[10]), .Y(n1491) );
  NAND2X1 U2708 ( .A(n711), .B(n714), .Y(n715) );
  NAND4X1 U2709 ( .A(n1633), .B(n1634), .C(n1635), .D(n1636), .Y(n714) );
  NOR4BX1 U2710 ( .AN(n711), .B(n1637), .C(n1638), .D(n1639), .Y(n1636) );
  XOR2X1 U2711 ( .A(\iforward/BUS937[0] ), .B(BUS18211[0]), .Y(n1639) );
  XOR2X1 U2712 ( .A(\iforward/BUS937[1] ), .B(BUS18211[1]), .Y(n1638) );
  XOR2X1 U2713 ( .A(\iforward/BUS937[3] ), .B(n1640), .Y(n1635) );
  XOR2X1 U2714 ( .A(\iforward/BUS937[4] ), .B(n1641), .Y(n1634) );
  XOR2X1 U2715 ( .A(\iforward/BUS937[2] ), .B(n1642), .Y(n1633) );
  NAND4X1 U2716 ( .A(n1643), .B(n1572), .C(n1644), .D(n1645), .Y(n711) );
  NOR3X1 U2717 ( .A(n1646), .B(n1647), .C(n1648), .Y(n1645) );
  XOR2X1 U2718 ( .A(\iforward/BUS937[2] ), .B(BUS1724[2]), .Y(n1648) );
  XOR2X1 U2719 ( .A(\iforward/BUS937[4] ), .B(BUS1724[4]), .Y(n1647) );
  XOR2X1 U2720 ( .A(\iforward/BUS937[3] ), .B(BUS1724[3]), .Y(n1646) );
  XOR2X1 U2721 ( .A(\iforward/BUS937[0] ), .B(n1578), .Y(n1644) );
  XOR2X1 U2722 ( .A(\iforward/BUS937[1] ), .B(n1579), .Y(n1643) );
  OAI221X1 U2723 ( .A0(n314), .A1(n299), .B0(n320), .B1(n300), .C0(n1649), .Y(
        BUS775[4]) );
  OAI221X1 U2724 ( .A0(n313), .A1(n299), .B0(n319), .B1(n300), .C0(n1649), .Y(
        BUS775[3]) );
  OAI221X1 U2725 ( .A0(n312), .A1(n299), .B0(n318), .B1(n300), .C0(n1649), .Y(
        BUS775[2]) );
  OAI221X1 U2726 ( .A0(n311), .A1(n299), .B0(n316), .B1(n300), .C0(n1649), .Y(
        BUS775[1]) );
  OAI221X1 U2727 ( .A0(n310), .A1(n299), .B0(n315), .B1(n300), .C0(n1649), .Y(
        BUS775[0]) );
  OR2X1 U2728 ( .A(n299), .B(n300), .Y(n1649) );
  OAI22X1 U2729 ( .A0(n308), .A1(n1650), .B0(n332), .B1(n1651), .Y(BUS7219[9])
         );
  OAI22X1 U2730 ( .A0(n307), .A1(n1650), .B0(n331), .B1(n1651), .Y(BUS7219[8])
         );
  OAI22X1 U2731 ( .A0(n332), .A1(n1650), .B0(n330), .B1(n1651), .Y(BUS7219[7])
         );
  OAI22X1 U2732 ( .A0(n331), .A1(n1650), .B0(n329), .B1(n1651), .Y(BUS7219[6])
         );
  OAI22X1 U2733 ( .A0(n330), .A1(n1650), .B0(n328), .B1(n1651), .Y(BUS7219[5])
         );
  OAI222X1 U2734 ( .A0(n309), .A1(n1652), .B0(n327), .B1(n1651), .C0(n329), 
        .C1(n1650), .Y(BUS7219[4]) );
  OAI222X1 U2735 ( .A0(n308), .A1(n1652), .B0(n326), .B1(n1651), .C0(n328), 
        .C1(n1650), .Y(BUS7219[3]) );
  OAI21X1 U2736 ( .A0(n314), .A1(n1653), .B0(n1654), .Y(BUS7219[31]) );
  OAI21X1 U2737 ( .A0(n313), .A1(n1653), .B0(n1654), .Y(BUS7219[30]) );
  OAI222X1 U2738 ( .A0(n307), .A1(n1652), .B0(n317), .B1(n1651), .C0(n327), 
        .C1(n1650), .Y(BUS7219[2]) );
  OAI21X1 U2739 ( .A0(n312), .A1(n1653), .B0(n1654), .Y(BUS7219[29]) );
  OAI21X1 U2740 ( .A0(n311), .A1(n1653), .B0(n1654), .Y(BUS7219[28]) );
  OAI221X1 U2741 ( .A0(n310), .A1(n1653), .B0(n325), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[27]) );
  OAI221X1 U2742 ( .A0(n309), .A1(n1653), .B0(n324), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[26]) );
  OAI221X1 U2743 ( .A0(n308), .A1(n1653), .B0(n323), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[25]) );
  OAI221X1 U2744 ( .A0(n307), .A1(n1653), .B0(n322), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[24]) );
  OAI221X1 U2745 ( .A0(n332), .A1(n1653), .B0(n321), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[23]) );
  OAI221X1 U2746 ( .A0(n331), .A1(n1653), .B0(n320), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[22]) );
  OAI221X1 U2747 ( .A0(n330), .A1(n1653), .B0(n319), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[21]) );
  OAI221X1 U2748 ( .A0(n329), .A1(n1653), .B0(n318), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[20]) );
  OAI22X1 U2749 ( .A0(n326), .A1(n1650), .B0(n332), .B1(n1652), .Y(BUS7219[1])
         );
  OAI221X1 U2750 ( .A0(n328), .A1(n1653), .B0(n316), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[19]) );
  OAI221X1 U2751 ( .A0(n327), .A1(n1653), .B0(n315), .B1(n1655), .C0(n1654), 
        .Y(BUS7219[18]) );
  OAI2BB1X1 U2752 ( .A0N(n1656), .A1N(n1657), .B0(n44), .Y(n1654) );
  CLKINVX1 U2753 ( .A(n1658), .Y(n1655) );
  OAI2BB2X1 U2754 ( .B0(n326), .B1(n1653), .A0N(n44), .A1N(n1659), .Y(
        BUS7219[17]) );
  OAI21X1 U2755 ( .A0(n42), .A1(n296), .B0(n1656), .Y(n1659) );
  OAI222X1 U2756 ( .A0(n313), .A1(n1651), .B0(n317), .B1(n1653), .C0(n314), 
        .C1(n1657), .Y(BUS7219[16]) );
  OR2X1 U2757 ( .A(n298), .B(n297), .Y(n1653) );
  OAI22X1 U2758 ( .A0(n314), .A1(n1650), .B0(n312), .B1(n1651), .Y(BUS7219[15]) );
  OAI22X1 U2759 ( .A0(n313), .A1(n1650), .B0(n311), .B1(n1651), .Y(BUS7219[14]) );
  OAI22X1 U2760 ( .A0(n312), .A1(n1650), .B0(n310), .B1(n1651), .Y(BUS7219[13]) );
  OAI22X1 U2761 ( .A0(n311), .A1(n1650), .B0(n309), .B1(n1651), .Y(BUS7219[12]) );
  OAI22X1 U2762 ( .A0(n310), .A1(n1650), .B0(n308), .B1(n1651), .Y(BUS7219[11]) );
  OAI22X1 U2763 ( .A0(n309), .A1(n1650), .B0(n307), .B1(n1651), .Y(BUS7219[10]) );
  AOI2BB1X1 U2764 ( .A0N(n298), .A1N(n1656), .B0(n1658), .Y(n1651) );
  NOR3X1 U2765 ( .A(n296), .B(n297), .C(n42), .Y(n1658) );
  NAND2X1 U2766 ( .A(n297), .B(n296), .Y(n1656) );
  OAI22X1 U2767 ( .A0(n317), .A1(n1650), .B0(n331), .B1(n1652), .Y(BUS7219[0])
         );
  OR2X1 U2768 ( .A(n298), .B(n296), .Y(n1652) );
  CLKINVX1 U2769 ( .A(n1660), .Y(n1650) );
  OAI2BB1X1 U2770 ( .A0N(n296), .A1N(n298), .B0(n1657), .Y(n1660) );
  NAND2X1 U2771 ( .A(n297), .B(n298), .Y(n1657) );
  OAI221X1 U2772 ( .A0(n1585), .A1(n1661), .B0(n1586), .B1(n1662), .C0(n1663), 
        .Y(BUS7160[9]) );
  AOI22X1 U2773 ( .A0(\iRF_stage/reg_bank/N1111 ), .A1(n1664), .B0(n1665), 
        .B1(n3), .Y(n1663) );
  OAI221X1 U2774 ( .A0(n1587), .A1(n1661), .B0(n1588), .B1(n1662), .C0(n1666), 
        .Y(BUS7160[8]) );
  AOI22X1 U2775 ( .A0(\iRF_stage/reg_bank/N1112 ), .A1(n1664), .B0(n1665), 
        .B1(n4), .Y(n1666) );
  OAI221X1 U2776 ( .A0(n718), .A1(n1661), .B0(n719), .B1(n1662), .C0(n1667), 
        .Y(BUS7160[7]) );
  AOI22X1 U2777 ( .A0(\iRF_stage/reg_bank/N1113 ), .A1(n1664), .B0(n1665), 
        .B1(n5), .Y(n1667) );
  OAI221X1 U2778 ( .A0(n721), .A1(n1661), .B0(n722), .B1(n1662), .C0(n1668), 
        .Y(BUS7160[6]) );
  AOI22X1 U2779 ( .A0(\iRF_stage/reg_bank/N1114 ), .A1(n1664), .B0(n1665), 
        .B1(n6), .Y(n1668) );
  OAI221X1 U2780 ( .A0(n724), .A1(n1661), .B0(n725), .B1(n1662), .C0(n1669), 
        .Y(BUS7160[5]) );
  AOI22X1 U2781 ( .A0(\iRF_stage/reg_bank/N1115 ), .A1(n1664), .B0(n1665), 
        .B1(n7), .Y(n1669) );
  OAI221X1 U2782 ( .A0(n727), .A1(n1661), .B0(n728), .B1(n1662), .C0(n1670), 
        .Y(BUS7160[4]) );
  AOI22X1 U2783 ( .A0(\iRF_stage/reg_bank/N1116 ), .A1(n1664), .B0(n1665), 
        .B1(n8), .Y(n1670) );
  OAI221X1 U2784 ( .A0(n730), .A1(n1661), .B0(n731), .B1(n1662), .C0(n1671), 
        .Y(BUS7160[3]) );
  AOI22X1 U2785 ( .A0(\iRF_stage/reg_bank/N1117 ), .A1(n1664), .B0(n1665), 
        .B1(n9), .Y(n1671) );
  OAI221X1 U2786 ( .A0(n1589), .A1(n1661), .B0(n1590), .B1(n1662), .C0(n1672), 
        .Y(BUS7160[31]) );
  AOI22X1 U2787 ( .A0(\iRF_stage/reg_bank/N1089 ), .A1(n1664), .B0(n1665), 
        .B1(n10), .Y(n1672) );
  OAI221X1 U2788 ( .A0(n1591), .A1(n1661), .B0(n1592), .B1(n1662), .C0(n1673), 
        .Y(BUS7160[30]) );
  AOI22X1 U2789 ( .A0(\iRF_stage/reg_bank/N1090 ), .A1(n1664), .B0(n1665), 
        .B1(n11), .Y(n1673) );
  OAI221X1 U2790 ( .A0(n733), .A1(n1661), .B0(n734), .B1(n1662), .C0(n1674), 
        .Y(BUS7160[2]) );
  AOI22X1 U2791 ( .A0(\iRF_stage/reg_bank/N1118 ), .A1(n1664), .B0(n1665), 
        .B1(n12), .Y(n1674) );
  OAI221X1 U2792 ( .A0(n1593), .A1(n1661), .B0(n1594), .B1(n1662), .C0(n1675), 
        .Y(BUS7160[29]) );
  AOI22X1 U2793 ( .A0(\iRF_stage/reg_bank/N1091 ), .A1(n1664), .B0(n1665), 
        .B1(n13), .Y(n1675) );
  OAI221X1 U2794 ( .A0(n1595), .A1(n1661), .B0(n1596), .B1(n1662), .C0(n1676), 
        .Y(BUS7160[28]) );
  AOI22X1 U2795 ( .A0(\iRF_stage/reg_bank/N1092 ), .A1(n1664), .B0(n1665), 
        .B1(n14), .Y(n1676) );
  OAI221X1 U2796 ( .A0(n1597), .A1(n1661), .B0(n1598), .B1(n1662), .C0(n1677), 
        .Y(BUS7160[27]) );
  AOI22X1 U2797 ( .A0(\iRF_stage/reg_bank/N1093 ), .A1(n1664), .B0(n1665), 
        .B1(n15), .Y(n1677) );
  OAI221X1 U2798 ( .A0(n1599), .A1(n1661), .B0(n1600), .B1(n1662), .C0(n1678), 
        .Y(BUS7160[26]) );
  AOI22X1 U2799 ( .A0(\iRF_stage/reg_bank/N1094 ), .A1(n1664), .B0(n1665), 
        .B1(n16), .Y(n1678) );
  OAI221X1 U2800 ( .A0(n1601), .A1(n1661), .B0(n1602), .B1(n1662), .C0(n1679), 
        .Y(BUS7160[25]) );
  AOI22X1 U2801 ( .A0(\iRF_stage/reg_bank/N1095 ), .A1(n1664), .B0(n1665), 
        .B1(n17), .Y(n1679) );
  OAI221X1 U2802 ( .A0(n1603), .A1(n1661), .B0(n1604), .B1(n1662), .C0(n1680), 
        .Y(BUS7160[24]) );
  AOI22X1 U2803 ( .A0(\iRF_stage/reg_bank/N1096 ), .A1(n1664), .B0(n1665), 
        .B1(n18), .Y(n1680) );
  OAI221X1 U2804 ( .A0(n1605), .A1(n1661), .B0(n1606), .B1(n1662), .C0(n1681), 
        .Y(BUS7160[23]) );
  AOI22X1 U2805 ( .A0(\iRF_stage/reg_bank/N1097 ), .A1(n1664), .B0(n1665), 
        .B1(n19), .Y(n1681) );
  OAI221X1 U2806 ( .A0(n1607), .A1(n1661), .B0(n1608), .B1(n1662), .C0(n1682), 
        .Y(BUS7160[22]) );
  AOI22X1 U2807 ( .A0(\iRF_stage/reg_bank/N1098 ), .A1(n1664), .B0(n1665), 
        .B1(n20), .Y(n1682) );
  OAI221X1 U2808 ( .A0(n1609), .A1(n1661), .B0(n1610), .B1(n1662), .C0(n1683), 
        .Y(BUS7160[21]) );
  AOI22X1 U2809 ( .A0(\iRF_stage/reg_bank/N1099 ), .A1(n1664), .B0(n1665), 
        .B1(n21), .Y(n1683) );
  OAI221X1 U2810 ( .A0(n1611), .A1(n1661), .B0(n1612), .B1(n1662), .C0(n1684), 
        .Y(BUS7160[20]) );
  AOI22X1 U2811 ( .A0(\iRF_stage/reg_bank/N1100 ), .A1(n1664), .B0(n1665), 
        .B1(n22), .Y(n1684) );
  OAI221X1 U2812 ( .A0(n712), .A1(n1661), .B0(n713), .B1(n1662), .C0(n1685), 
        .Y(BUS7160[1]) );
  AOI22X1 U2813 ( .A0(\iRF_stage/reg_bank/N1119 ), .A1(n1664), .B0(n1665), 
        .B1(n23), .Y(n1685) );
  OAI221X1 U2814 ( .A0(n1613), .A1(n1661), .B0(n1614), .B1(n1662), .C0(n1686), 
        .Y(BUS7160[19]) );
  AOI22X1 U2815 ( .A0(\iRF_stage/reg_bank/N1101 ), .A1(n1664), .B0(n1665), 
        .B1(n24), .Y(n1686) );
  OAI221X1 U2816 ( .A0(n1615), .A1(n1661), .B0(n1616), .B1(n1662), .C0(n1687), 
        .Y(BUS7160[18]) );
  AOI22X1 U2817 ( .A0(\iRF_stage/reg_bank/N1102 ), .A1(n1664), .B0(n1665), 
        .B1(n25), .Y(n1687) );
  OAI221X1 U2818 ( .A0(n1617), .A1(n1661), .B0(n1618), .B1(n1662), .C0(n1688), 
        .Y(BUS7160[17]) );
  AOI22X1 U2819 ( .A0(\iRF_stage/reg_bank/N1103 ), .A1(n1664), .B0(n1665), 
        .B1(n26), .Y(n1688) );
  OAI221X1 U2820 ( .A0(n1619), .A1(n1661), .B0(n1620), .B1(n1662), .C0(n1689), 
        .Y(BUS7160[16]) );
  AOI22X1 U2821 ( .A0(\iRF_stage/reg_bank/N1104 ), .A1(n1664), .B0(n1665), 
        .B1(n27), .Y(n1689) );
  OAI221X1 U2822 ( .A0(n1621), .A1(n1661), .B0(n1622), .B1(n1662), .C0(n1690), 
        .Y(BUS7160[15]) );
  AOI22X1 U2823 ( .A0(\iRF_stage/reg_bank/N1105 ), .A1(n1664), .B0(n1665), 
        .B1(n28), .Y(n1690) );
  OAI221X1 U2824 ( .A0(n1623), .A1(n1661), .B0(n1624), .B1(n1662), .C0(n1691), 
        .Y(BUS7160[14]) );
  AOI22X1 U2825 ( .A0(\iRF_stage/reg_bank/N1106 ), .A1(n1664), .B0(n1665), 
        .B1(n29), .Y(n1691) );
  OAI221X1 U2826 ( .A0(n1625), .A1(n1661), .B0(n1626), .B1(n1662), .C0(n1692), 
        .Y(BUS7160[13]) );
  AOI22X1 U2827 ( .A0(\iRF_stage/reg_bank/N1107 ), .A1(n1664), .B0(n1665), 
        .B1(n30), .Y(n1692) );
  OAI221X1 U2828 ( .A0(n1627), .A1(n1661), .B0(n1628), .B1(n1662), .C0(n1693), 
        .Y(BUS7160[12]) );
  AOI22X1 U2829 ( .A0(\iRF_stage/reg_bank/N1108 ), .A1(n1664), .B0(n1665), 
        .B1(n31), .Y(n1693) );
  OAI221X1 U2830 ( .A0(n1629), .A1(n1661), .B0(n1630), .B1(n1662), .C0(n1694), 
        .Y(BUS7160[11]) );
  AOI22X1 U2831 ( .A0(\iRF_stage/reg_bank/N1109 ), .A1(n1664), .B0(n1665), 
        .B1(n32), .Y(n1694) );
  OAI221X1 U2832 ( .A0(n1631), .A1(n1661), .B0(n1632), .B1(n1662), .C0(n1695), 
        .Y(BUS7160[10]) );
  AOI22X1 U2833 ( .A0(\iRF_stage/reg_bank/N1110 ), .A1(n1664), .B0(n1665), 
        .B1(n33), .Y(n1695) );
  OAI221X1 U2834 ( .A0(n736), .A1(n1661), .B0(n737), .B1(n1662), .C0(n1696), 
        .Y(BUS7160[0]) );
  AOI22X1 U2835 ( .A0(\iRF_stage/reg_bank/N1120 ), .A1(n1664), .B0(n1665), 
        .B1(n34), .Y(n1696) );
  AND3X2 U2836 ( .A(n1697), .B(n1698), .C(n1699), .Y(n1665) );
  CLKINVX1 U2837 ( .A(n1700), .Y(n1697) );
  AND3X2 U2838 ( .A(n1698), .B(n1699), .C(n1700), .Y(n1664) );
  NAND4X1 U2839 ( .A(n1701), .B(n1702), .C(\iRF_stage/reg_bank/r_wren ), .D(
        n1703), .Y(n1700) );
  NOR3X1 U2840 ( .A(n1704), .B(n1705), .C(n1706), .Y(n1703) );
  XOR2X1 U2841 ( .A(n333), .B(n630), .Y(n1706) );
  XOR2X1 U2842 ( .A(n339), .B(n642), .Y(n1705) );
  XOR2X1 U2843 ( .A(n342), .B(n620), .Y(n1704) );
  CLKINVX1 U2844 ( .A(\iRF_stage/reg_bank/r_wraddress[3] ), .Y(n620) );
  XOR2X1 U2845 ( .A(\iRF_stage/reg_bank/r_wraddress[1] ), .B(n340), .Y(n1702)
         );
  XOR2X1 U2846 ( .A(\iRF_stage/reg_bank/r_wraddress[2] ), .B(n341), .Y(n1701)
         );
  NAND4X1 U2847 ( .A(n342), .B(n341), .C(n1707), .D(n340), .Y(n1699) );
  AND2X1 U2848 ( .A(n333), .B(n339), .Y(n1707) );
  AND2X1 U2849 ( .A(n1661), .B(n1662), .Y(n1698) );
  NAND4X1 U2850 ( .A(n1708), .B(n1709), .C(n1563), .D(n1710), .Y(n1662) );
  NOR4BX1 U2851 ( .AN(n1661), .B(n1711), .C(n1712), .D(n1713), .Y(n1710) );
  XOR2X1 U2852 ( .A(n1641), .B(n320), .Y(n1713) );
  XOR2X1 U2853 ( .A(n1569), .B(n315), .Y(n1712) );
  XOR2X1 U2854 ( .A(n1570), .B(n316), .Y(n1711) );
  XOR2X1 U2855 ( .A(n318), .B(BUS18211[2]), .Y(n1709) );
  XOR2X1 U2856 ( .A(n319), .B(BUS18211[3]), .Y(n1708) );
  NAND4X1 U2857 ( .A(n1714), .B(n1715), .C(n1572), .D(n1716), .Y(n1661) );
  NOR3X1 U2858 ( .A(n1717), .B(n1718), .C(n1719), .Y(n1716) );
  XOR2X1 U2859 ( .A(n1578), .B(n315), .Y(n1719) );
  XOR2X1 U2860 ( .A(n1579), .B(n316), .Y(n1718) );
  XOR2X1 U2861 ( .A(n1720), .B(n320), .Y(n1717) );
  XOR2X1 U2862 ( .A(n318), .B(BUS1724[2]), .Y(n1715) );
  XOR2X1 U2863 ( .A(n319), .B(BUS1724[3]), .Y(n1714) );
  OAI221X1 U2864 ( .A0(n1585), .A1(n1721), .B0(n1586), .B1(n1722), .C0(n1723), 
        .Y(BUS24839[9]) );
  AOI22X1 U2865 ( .A0(\iRF_stage/reg_bank/N1074 ), .A1(n1724), .B0(n1725), 
        .B1(n3), .Y(n1723) );
  CLKINVX1 U2866 ( .A(cop_addr_o[9]), .Y(n1585) );
  OAI221X1 U2867 ( .A0(n1587), .A1(n1721), .B0(n1588), .B1(n1722), .C0(n1726), 
        .Y(BUS24839[8]) );
  AOI22X1 U2868 ( .A0(\iRF_stage/reg_bank/N1075 ), .A1(n1724), .B0(n1725), 
        .B1(n4), .Y(n1726) );
  CLKINVX1 U2869 ( .A(cop_addr_o[8]), .Y(n1587) );
  OAI221X1 U2870 ( .A0(n718), .A1(n1721), .B0(n719), .B1(n1722), .C0(n1727), 
        .Y(BUS24839[7]) );
  AOI22X1 U2871 ( .A0(\iRF_stage/reg_bank/N1076 ), .A1(n1724), .B0(n1725), 
        .B1(n5), .Y(n1727) );
  CLKINVX1 U2872 ( .A(cop_addr_o[7]), .Y(n718) );
  OAI221X1 U2873 ( .A0(n721), .A1(n1721), .B0(n722), .B1(n1722), .C0(n1728), 
        .Y(BUS24839[6]) );
  AOI22X1 U2874 ( .A0(\iRF_stage/reg_bank/N1077 ), .A1(n1724), .B0(n1725), 
        .B1(n6), .Y(n1728) );
  CLKINVX1 U2875 ( .A(cop_addr_o[6]), .Y(n721) );
  OAI221X1 U2876 ( .A0(n724), .A1(n1721), .B0(n725), .B1(n1722), .C0(n1729), 
        .Y(BUS24839[5]) );
  AOI22X1 U2877 ( .A0(\iRF_stage/reg_bank/N1078 ), .A1(n1724), .B0(n1725), 
        .B1(n7), .Y(n1729) );
  CLKINVX1 U2878 ( .A(cop_addr_o[5]), .Y(n724) );
  OAI221X1 U2879 ( .A0(n727), .A1(n1721), .B0(n728), .B1(n1722), .C0(n1730), 
        .Y(BUS24839[4]) );
  AOI22X1 U2880 ( .A0(\iRF_stage/reg_bank/N1079 ), .A1(n1724), .B0(n1725), 
        .B1(n8), .Y(n1730) );
  CLKINVX1 U2881 ( .A(cop_addr_o[4]), .Y(n727) );
  OAI221X1 U2882 ( .A0(n730), .A1(n1721), .B0(n731), .B1(n1722), .C0(n1731), 
        .Y(BUS24839[3]) );
  AOI22X1 U2883 ( .A0(\iRF_stage/reg_bank/N1080 ), .A1(n1724), .B0(n1725), 
        .B1(n9), .Y(n1731) );
  CLKINVX1 U2884 ( .A(cop_addr_o[3]), .Y(n730) );
  OAI221X1 U2885 ( .A0(n1589), .A1(n1721), .B0(n1590), .B1(n1722), .C0(n1732), 
        .Y(BUS24839[31]) );
  AOI22X1 U2886 ( .A0(\iRF_stage/reg_bank/N1052 ), .A1(n1724), .B0(n1725), 
        .B1(n10), .Y(n1732) );
  CLKINVX1 U2887 ( .A(cop_addr_o[31]), .Y(n1589) );
  OAI221X1 U2888 ( .A0(n1591), .A1(n1721), .B0(n1592), .B1(n1722), .C0(n1733), 
        .Y(BUS24839[30]) );
  AOI22X1 U2889 ( .A0(\iRF_stage/reg_bank/N1053 ), .A1(n1724), .B0(n1725), 
        .B1(n11), .Y(n1733) );
  CLKINVX1 U2890 ( .A(cop_addr_o[30]), .Y(n1591) );
  OAI221X1 U2891 ( .A0(n733), .A1(n1721), .B0(n734), .B1(n1722), .C0(n1734), 
        .Y(BUS24839[2]) );
  AOI22X1 U2892 ( .A0(\iRF_stage/reg_bank/N1081 ), .A1(n1724), .B0(n1725), 
        .B1(n12), .Y(n1734) );
  CLKINVX1 U2893 ( .A(cop_addr_o[2]), .Y(n733) );
  OAI221X1 U2894 ( .A0(n1593), .A1(n1721), .B0(n1594), .B1(n1722), .C0(n1735), 
        .Y(BUS24839[29]) );
  AOI22X1 U2895 ( .A0(\iRF_stage/reg_bank/N1054 ), .A1(n1724), .B0(n1725), 
        .B1(n13), .Y(n1735) );
  CLKINVX1 U2896 ( .A(cop_addr_o[29]), .Y(n1593) );
  OAI221X1 U2897 ( .A0(n1595), .A1(n1721), .B0(n1596), .B1(n1722), .C0(n1736), 
        .Y(BUS24839[28]) );
  AOI22X1 U2898 ( .A0(\iRF_stage/reg_bank/N1055 ), .A1(n1724), .B0(n1725), 
        .B1(n14), .Y(n1736) );
  CLKINVX1 U2899 ( .A(cop_addr_o[28]), .Y(n1595) );
  OAI221X1 U2900 ( .A0(n1597), .A1(n1721), .B0(n1598), .B1(n1722), .C0(n1737), 
        .Y(BUS24839[27]) );
  AOI22X1 U2901 ( .A0(\iRF_stage/reg_bank/N1056 ), .A1(n1724), .B0(n1725), 
        .B1(n15), .Y(n1737) );
  CLKINVX1 U2902 ( .A(cop_addr_o[27]), .Y(n1597) );
  OAI221X1 U2903 ( .A0(n1599), .A1(n1721), .B0(n1600), .B1(n1722), .C0(n1738), 
        .Y(BUS24839[26]) );
  AOI22X1 U2904 ( .A0(\iRF_stage/reg_bank/N1057 ), .A1(n1724), .B0(n1725), 
        .B1(n16), .Y(n1738) );
  CLKINVX1 U2905 ( .A(cop_addr_o[26]), .Y(n1599) );
  OAI221X1 U2906 ( .A0(n1601), .A1(n1721), .B0(n1602), .B1(n1722), .C0(n1739), 
        .Y(BUS24839[25]) );
  AOI22X1 U2907 ( .A0(\iRF_stage/reg_bank/N1058 ), .A1(n1724), .B0(n1725), 
        .B1(n17), .Y(n1739) );
  CLKINVX1 U2908 ( .A(cop_addr_o[25]), .Y(n1601) );
  OAI221X1 U2909 ( .A0(n1603), .A1(n1721), .B0(n1604), .B1(n1722), .C0(n1740), 
        .Y(BUS24839[24]) );
  AOI22X1 U2910 ( .A0(\iRF_stage/reg_bank/N1059 ), .A1(n1724), .B0(n1725), 
        .B1(n18), .Y(n1740) );
  CLKINVX1 U2911 ( .A(cop_addr_o[24]), .Y(n1603) );
  OAI221X1 U2912 ( .A0(n1605), .A1(n1721), .B0(n1606), .B1(n1722), .C0(n1741), 
        .Y(BUS24839[23]) );
  AOI22X1 U2913 ( .A0(\iRF_stage/reg_bank/N1060 ), .A1(n1724), .B0(n1725), 
        .B1(n19), .Y(n1741) );
  CLKINVX1 U2914 ( .A(cop_addr_o[23]), .Y(n1605) );
  OAI221X1 U2915 ( .A0(n1607), .A1(n1721), .B0(n1608), .B1(n1722), .C0(n1742), 
        .Y(BUS24839[22]) );
  AOI22X1 U2916 ( .A0(\iRF_stage/reg_bank/N1061 ), .A1(n1724), .B0(n1725), 
        .B1(n20), .Y(n1742) );
  CLKINVX1 U2917 ( .A(cop_addr_o[22]), .Y(n1607) );
  OAI221X1 U2918 ( .A0(n1609), .A1(n1721), .B0(n1610), .B1(n1722), .C0(n1743), 
        .Y(BUS24839[21]) );
  AOI22X1 U2919 ( .A0(\iRF_stage/reg_bank/N1062 ), .A1(n1724), .B0(n1725), 
        .B1(n21), .Y(n1743) );
  CLKINVX1 U2920 ( .A(cop_addr_o[21]), .Y(n1609) );
  OAI221X1 U2921 ( .A0(n1611), .A1(n1721), .B0(n1612), .B1(n1722), .C0(n1744), 
        .Y(BUS24839[20]) );
  AOI22X1 U2922 ( .A0(\iRF_stage/reg_bank/N1063 ), .A1(n1724), .B0(n1725), 
        .B1(n22), .Y(n1744) );
  CLKINVX1 U2923 ( .A(cop_addr_o[20]), .Y(n1611) );
  OAI221X1 U2924 ( .A0(n712), .A1(n1721), .B0(n713), .B1(n1722), .C0(n1745), 
        .Y(BUS24839[1]) );
  AOI22X1 U2925 ( .A0(\iRF_stage/reg_bank/N1082 ), .A1(n1724), .B0(n1725), 
        .B1(n23), .Y(n1745) );
  CLKINVX1 U2926 ( .A(cop_addr_o[1]), .Y(n712) );
  OAI221X1 U2927 ( .A0(n1613), .A1(n1721), .B0(n1614), .B1(n1722), .C0(n1746), 
        .Y(BUS24839[19]) );
  AOI22X1 U2928 ( .A0(\iRF_stage/reg_bank/N1064 ), .A1(n1724), .B0(n1725), 
        .B1(n24), .Y(n1746) );
  CLKINVX1 U2929 ( .A(cop_addr_o[19]), .Y(n1613) );
  OAI221X1 U2930 ( .A0(n1615), .A1(n1721), .B0(n1616), .B1(n1722), .C0(n1747), 
        .Y(BUS24839[18]) );
  AOI22X1 U2931 ( .A0(\iRF_stage/reg_bank/N1065 ), .A1(n1724), .B0(n1725), 
        .B1(n25), .Y(n1747) );
  CLKINVX1 U2932 ( .A(cop_addr_o[18]), .Y(n1615) );
  OAI221X1 U2933 ( .A0(n1617), .A1(n1721), .B0(n1618), .B1(n1722), .C0(n1748), 
        .Y(BUS24839[17]) );
  AOI22X1 U2934 ( .A0(\iRF_stage/reg_bank/N1066 ), .A1(n1724), .B0(n1725), 
        .B1(n26), .Y(n1748) );
  CLKINVX1 U2935 ( .A(cop_addr_o[17]), .Y(n1617) );
  OAI221X1 U2936 ( .A0(n1619), .A1(n1721), .B0(n1620), .B1(n1722), .C0(n1749), 
        .Y(BUS24839[16]) );
  AOI22X1 U2937 ( .A0(\iRF_stage/reg_bank/N1067 ), .A1(n1724), .B0(n1725), 
        .B1(n27), .Y(n1749) );
  CLKINVX1 U2938 ( .A(cop_addr_o[16]), .Y(n1619) );
  OAI221X1 U2939 ( .A0(n1621), .A1(n1721), .B0(n1622), .B1(n1722), .C0(n1750), 
        .Y(BUS24839[15]) );
  AOI22X1 U2940 ( .A0(\iRF_stage/reg_bank/N1068 ), .A1(n1724), .B0(n1725), 
        .B1(n28), .Y(n1750) );
  CLKINVX1 U2941 ( .A(cop_addr_o[15]), .Y(n1621) );
  OAI221X1 U2942 ( .A0(n1623), .A1(n1721), .B0(n1624), .B1(n1722), .C0(n1751), 
        .Y(BUS24839[14]) );
  AOI22X1 U2943 ( .A0(\iRF_stage/reg_bank/N1069 ), .A1(n1724), .B0(n1725), 
        .B1(n29), .Y(n1751) );
  CLKINVX1 U2944 ( .A(cop_addr_o[14]), .Y(n1623) );
  OAI221X1 U2945 ( .A0(n1625), .A1(n1721), .B0(n1626), .B1(n1722), .C0(n1752), 
        .Y(BUS24839[13]) );
  AOI22X1 U2946 ( .A0(\iRF_stage/reg_bank/N1070 ), .A1(n1724), .B0(n1725), 
        .B1(n30), .Y(n1752) );
  CLKINVX1 U2947 ( .A(cop_addr_o[13]), .Y(n1625) );
  OAI221X1 U2948 ( .A0(n1627), .A1(n1721), .B0(n1628), .B1(n1722), .C0(n1753), 
        .Y(BUS24839[12]) );
  AOI22X1 U2949 ( .A0(\iRF_stage/reg_bank/N1071 ), .A1(n1724), .B0(n1725), 
        .B1(n31), .Y(n1753) );
  CLKINVX1 U2950 ( .A(cop_addr_o[12]), .Y(n1627) );
  OAI221X1 U2951 ( .A0(n1629), .A1(n1721), .B0(n1630), .B1(n1722), .C0(n1754), 
        .Y(BUS24839[11]) );
  AOI22X1 U2952 ( .A0(\iRF_stage/reg_bank/N1072 ), .A1(n1724), .B0(n1725), 
        .B1(n32), .Y(n1754) );
  CLKINVX1 U2953 ( .A(cop_addr_o[11]), .Y(n1629) );
  OAI221X1 U2954 ( .A0(n1631), .A1(n1721), .B0(n1632), .B1(n1722), .C0(n1755), 
        .Y(BUS24839[10]) );
  AOI22X1 U2955 ( .A0(\iRF_stage/reg_bank/N1073 ), .A1(n1724), .B0(n1725), 
        .B1(n33), .Y(n1755) );
  CLKINVX1 U2956 ( .A(cop_addr_o[10]), .Y(n1631) );
  OAI221X1 U2957 ( .A0(n736), .A1(n1721), .B0(n737), .B1(n1722), .C0(n1756), 
        .Y(BUS24839[0]) );
  AOI22X1 U2958 ( .A0(\iRF_stage/reg_bank/N1083 ), .A1(n1724), .B0(n1725), 
        .B1(n34), .Y(n1756) );
  AND3X2 U2959 ( .A(n1757), .B(n1758), .C(n1759), .Y(n1725) );
  CLKINVX1 U2960 ( .A(n1760), .Y(n1757) );
  AND3X2 U2961 ( .A(n1758), .B(n1759), .C(n1760), .Y(n1724) );
  NAND4X1 U2962 ( .A(n1761), .B(n1762), .C(\iRF_stage/reg_bank/r_wren ), .D(
        n1763), .Y(n1760) );
  NOR3X1 U2963 ( .A(n1764), .B(n1765), .C(n1766), .Y(n1763) );
  XOR2X1 U2964 ( .A(n334), .B(n642), .Y(n1766) );
  CLKINVX1 U2965 ( .A(\iRF_stage/reg_bank/r_wraddress[0] ), .Y(n642) );
  XOR2X1 U2966 ( .A(n335), .B(n639), .Y(n1765) );
  CLKINVX1 U2967 ( .A(\iRF_stage/reg_bank/r_wraddress[1] ), .Y(n639) );
  XOR2X1 U2968 ( .A(n338), .B(n630), .Y(n1764) );
  CLKINVX1 U2969 ( .A(\iRF_stage/reg_bank/r_wraddress[4] ), .Y(n630) );
  XOR2X1 U2970 ( .A(\iRF_stage/reg_bank/r_wraddress[2] ), .B(n336), .Y(n1762)
         );
  XOR2X1 U2971 ( .A(\iRF_stage/reg_bank/r_wraddress[3] ), .B(n337), .Y(n1761)
         );
  NAND4X1 U2972 ( .A(n338), .B(n337), .C(n1767), .D(n336), .Y(n1759) );
  AND2X1 U2973 ( .A(n334), .B(n335), .Y(n1767) );
  AND2X1 U2974 ( .A(n1721), .B(n1722), .Y(n1758) );
  NAND4X1 U2975 ( .A(n1768), .B(n1769), .C(n1563), .D(n1770), .Y(n1722) );
  NOR4BX1 U2976 ( .AN(n1721), .B(n1771), .C(n1772), .D(n1773), .Y(n1770) );
  XOR2X1 U2977 ( .A(n325), .B(n1641), .Y(n1773) );
  XOR2X1 U2978 ( .A(n321), .B(n1569), .Y(n1772) );
  CLKINVX1 U2979 ( .A(BUS18211[0]), .Y(n1569) );
  XOR2X1 U2980 ( .A(n322), .B(n1570), .Y(n1771) );
  CLKINVX1 U2981 ( .A(BUS18211[1]), .Y(n1570) );
  CLKINVX1 U2982 ( .A(n1637), .Y(n1563) );
  OAI31X1 U2983 ( .A0(n1774), .A1(BUS18211[1]), .A2(BUS18211[0]), .B0(NET1375), 
        .Y(n1637) );
  NAND3X1 U2984 ( .A(n1640), .B(n1641), .C(n1642), .Y(n1774) );
  CLKINVX1 U2985 ( .A(BUS18211[2]), .Y(n1642) );
  CLKINVX1 U2986 ( .A(BUS18211[4]), .Y(n1641) );
  CLKINVX1 U2987 ( .A(BUS18211[3]), .Y(n1640) );
  XOR2X1 U2988 ( .A(n323), .B(BUS18211[2]), .Y(n1769) );
  XOR2X1 U2989 ( .A(n324), .B(BUS18211[3]), .Y(n1768) );
  NAND4X1 U2990 ( .A(n1775), .B(n1776), .C(n1572), .D(n1777), .Y(n1721) );
  NOR3X1 U2991 ( .A(n1778), .B(n1779), .C(n1780), .Y(n1777) );
  XOR2X1 U2992 ( .A(n321), .B(n1578), .Y(n1780) );
  CLKINVX1 U2993 ( .A(BUS1724[0]), .Y(n1578) );
  XOR2X1 U2994 ( .A(n322), .B(n1579), .Y(n1779) );
  CLKINVX1 U2995 ( .A(BUS1724[1]), .Y(n1579) );
  XOR2X1 U2996 ( .A(n325), .B(n1720), .Y(n1778) );
  CLKINVX1 U2997 ( .A(BUS1724[4]), .Y(n1720) );
  CLKINVX1 U2998 ( .A(n1781), .Y(n1572) );
  OAI31X1 U2999 ( .A0(n1782), .A1(BUS1724[1]), .A2(BUS1724[0]), .B0(NET767), 
        .Y(n1781) );
  OR3X1 U3000 ( .A(BUS1724[3]), .B(BUS1724[4]), .C(BUS1724[2]), .Y(n1782) );
  XOR2X1 U3001 ( .A(n323), .B(BUS1724[2]), .Y(n1776) );
  XOR2X1 U3002 ( .A(n324), .B(BUS1724[3]), .Y(n1775) );
  CLKINVX1 U3003 ( .A(cop_addr_o[0]), .Y(n736) );
  NOR2X1 U3004 ( .A(n1783), .B(n35), .Y(BUS22401[9]) );
  AOI221XL U3005 ( .A0(din[25]), .A1(n1784), .B0(din[9]), .B1(n1785), .C0(
        n1786), .Y(n1783) );
  NOR2X1 U3006 ( .A(n1787), .B(n35), .Y(BUS22401[8]) );
  AOI221XL U3007 ( .A0(din[24]), .A1(n1784), .B0(din[8]), .B1(n1785), .C0(
        n1786), .Y(n1787) );
  NOR2X1 U3008 ( .A(n1788), .B(n35), .Y(BUS22401[7]) );
  AOI222XL U3009 ( .A0(din[23]), .A1(n1789), .B0(n1790), .B1(n1791), .C0(
        din[7]), .C1(n1792), .Y(n1788) );
  NOR2X1 U3010 ( .A(\MEM_CTL/BUS629[0] ), .B(n1793), .Y(n1790) );
  NOR2X1 U3011 ( .A(n1794), .B(n35), .Y(BUS22401[6]) );
  AOI221XL U3012 ( .A0(din[6]), .A1(n1792), .B0(din[22]), .B1(n1789), .C0(
        n1795), .Y(n1794) );
  OAI22X1 U3013 ( .A0(n1796), .A1(n1797), .B0(n1798), .B1(n1799), .Y(n1795) );
  CLKINVX1 U3014 ( .A(din[14]), .Y(n1799) );
  CLKINVX1 U3015 ( .A(din[30]), .Y(n1797) );
  NOR2X1 U3016 ( .A(n1800), .B(n35), .Y(BUS22401[5]) );
  AOI221XL U3017 ( .A0(din[5]), .A1(n1792), .B0(din[21]), .B1(n1789), .C0(
        n1801), .Y(n1800) );
  OAI22X1 U3018 ( .A0(n1796), .A1(n1802), .B0(n1798), .B1(n1803), .Y(n1801) );
  CLKINVX1 U3019 ( .A(din[13]), .Y(n1803) );
  CLKINVX1 U3020 ( .A(din[29]), .Y(n1802) );
  NOR2X1 U3021 ( .A(n1804), .B(n35), .Y(BUS22401[4]) );
  AOI221XL U3022 ( .A0(din[4]), .A1(n1792), .B0(din[20]), .B1(n1789), .C0(
        n1805), .Y(n1804) );
  OAI22X1 U3023 ( .A0(n1796), .A1(n1806), .B0(n1798), .B1(n1807), .Y(n1805) );
  CLKINVX1 U3024 ( .A(din[12]), .Y(n1807) );
  CLKINVX1 U3025 ( .A(din[28]), .Y(n1806) );
  NOR2X1 U3026 ( .A(n1808), .B(n35), .Y(BUS22401[3]) );
  AOI221XL U3027 ( .A0(din[3]), .A1(n1792), .B0(din[19]), .B1(n1789), .C0(
        n1809), .Y(n1808) );
  OAI22X1 U3028 ( .A0(n1796), .A1(n1810), .B0(n1798), .B1(n1811), .Y(n1809) );
  CLKINVX1 U3029 ( .A(din[11]), .Y(n1811) );
  CLKINVX1 U3030 ( .A(din[27]), .Y(n1810) );
  OAI2BB1X1 U3031 ( .A0N(n1812), .A1N(din[31]), .B0(n1813), .Y(BUS22401[31])
         );
  OAI2BB1X1 U3032 ( .A0N(din[30]), .A1N(n1812), .B0(n1813), .Y(BUS22401[30])
         );
  NOR2X1 U3033 ( .A(n1814), .B(n35), .Y(BUS22401[2]) );
  AOI221XL U3034 ( .A0(din[2]), .A1(n1792), .B0(din[18]), .B1(n1789), .C0(
        n1815), .Y(n1814) );
  OAI22X1 U3035 ( .A0(n1796), .A1(n1816), .B0(n1798), .B1(n1817), .Y(n1815) );
  CLKINVX1 U3036 ( .A(din[10]), .Y(n1817) );
  CLKINVX1 U3037 ( .A(din[26]), .Y(n1816) );
  OAI2BB1X1 U3038 ( .A0N(din[29]), .A1N(n1812), .B0(n1813), .Y(BUS22401[29])
         );
  OAI2BB1X1 U3039 ( .A0N(din[28]), .A1N(n1812), .B0(n1813), .Y(BUS22401[28])
         );
  OAI2BB1X1 U3040 ( .A0N(din[27]), .A1N(n1812), .B0(n1813), .Y(BUS22401[27])
         );
  OAI2BB1X1 U3041 ( .A0N(n1812), .A1N(din[26]), .B0(n1813), .Y(BUS22401[26])
         );
  OAI2BB1X1 U3042 ( .A0N(din[25]), .A1N(n1812), .B0(n1813), .Y(BUS22401[25])
         );
  OAI2BB1X1 U3043 ( .A0N(din[24]), .A1N(n1812), .B0(n1813), .Y(BUS22401[24])
         );
  OAI2BB1X1 U3044 ( .A0N(din[23]), .A1N(n1812), .B0(n1813), .Y(BUS22401[23])
         );
  OAI2BB1X1 U3045 ( .A0N(din[22]), .A1N(n1812), .B0(n1813), .Y(BUS22401[22])
         );
  OAI2BB1X1 U3046 ( .A0N(din[21]), .A1N(n1812), .B0(n1813), .Y(BUS22401[21])
         );
  OAI2BB1X1 U3047 ( .A0N(din[20]), .A1N(n1812), .B0(n1813), .Y(BUS22401[20])
         );
  NOR2X1 U3048 ( .A(n1818), .B(n35), .Y(BUS22401[1]) );
  AOI221XL U3049 ( .A0(din[1]), .A1(n1792), .B0(din[17]), .B1(n1789), .C0(
        n1819), .Y(n1818) );
  OAI22X1 U3050 ( .A0(n1820), .A1(n1796), .B0(n1821), .B1(n1798), .Y(n1819) );
  CLKINVX1 U3051 ( .A(din[9]), .Y(n1821) );
  CLKINVX1 U3052 ( .A(din[25]), .Y(n1820) );
  OAI2BB1X1 U3053 ( .A0N(din[19]), .A1N(n1812), .B0(n1813), .Y(BUS22401[19])
         );
  OAI2BB1X1 U3054 ( .A0N(n1812), .A1N(din[18]), .B0(n1813), .Y(BUS22401[18])
         );
  OAI2BB1X1 U3055 ( .A0N(n1812), .A1N(din[17]), .B0(n1813), .Y(BUS22401[17])
         );
  OAI2BB1X1 U3056 ( .A0N(n1812), .A1N(din[16]), .B0(n1813), .Y(BUS22401[16])
         );
  CLKINVX1 U3057 ( .A(n1822), .Y(n1812) );
  OAI221X1 U3058 ( .A0(n1823), .A1(n1824), .B0(n1822), .B1(n1825), .C0(n1813), 
        .Y(BUS22401[15]) );
  OR2X1 U3059 ( .A(n35), .B(n1826), .Y(n1813) );
  AOI31X1 U3060 ( .A0(n1791), .A1(n1827), .A2(n277), .B0(n1786), .Y(n1826) );
  CLKINVX1 U3061 ( .A(n1823), .Y(n1791) );
  CLKINVX1 U3062 ( .A(din[15]), .Y(n1825) );
  NAND2X1 U3063 ( .A(n1828), .B(n276), .Y(n1822) );
  NAND2X1 U3064 ( .A(n276), .B(n1827), .Y(n1824) );
  NOR2X1 U3065 ( .A(n1829), .B(n35), .Y(BUS22401[14]) );
  AOI221XL U3066 ( .A0(din[30]), .A1(n1784), .B0(din[14]), .B1(n1785), .C0(
        n1786), .Y(n1829) );
  NOR2X1 U3067 ( .A(n1830), .B(n35), .Y(BUS22401[13]) );
  AOI221XL U3068 ( .A0(din[29]), .A1(n1784), .B0(din[13]), .B1(n1785), .C0(
        n1786), .Y(n1830) );
  NOR2X1 U3069 ( .A(n1831), .B(n35), .Y(BUS22401[12]) );
  AOI221XL U3070 ( .A0(din[28]), .A1(n1784), .B0(din[12]), .B1(n1785), .C0(
        n1786), .Y(n1831) );
  NOR2X1 U3071 ( .A(n1832), .B(n35), .Y(BUS22401[11]) );
  AOI221XL U3072 ( .A0(din[27]), .A1(n1784), .B0(din[11]), .B1(n1785), .C0(
        n1786), .Y(n1832) );
  NOR2X1 U3073 ( .A(n1833), .B(n35), .Y(BUS22401[10]) );
  AOI221XL U3074 ( .A0(din[26]), .A1(n1784), .B0(din[10]), .B1(n1785), .C0(
        n1786), .Y(n1833) );
  AND2X1 U3075 ( .A(n1834), .B(n1835), .Y(n1786) );
  MXI2X1 U3076 ( .A(n1823), .B(n1836), .S0(\MEM_CTL/BUS629[0] ), .Y(n1834) );
  MXI2X1 U3077 ( .A(din[23]), .B(din[7]), .S0(\MEM_CTL/BUS629[1] ), .Y(n1836)
         );
  MXI2X1 U3078 ( .A(din[31]), .B(din[15]), .S0(\MEM_CTL/BUS629[1] ), .Y(n1823)
         );
  CLKINVX1 U3079 ( .A(n1837), .Y(n1785) );
  CLKINVX1 U3080 ( .A(n1838), .Y(n1784) );
  NOR2X1 U3081 ( .A(n1839), .B(n35), .Y(BUS22401[0]) );
  AOI221XL U3082 ( .A0(din[0]), .A1(n1792), .B0(din[16]), .B1(n1789), .C0(
        n1840), .Y(n1839) );
  OAI22X1 U3083 ( .A0(n1841), .A1(n1796), .B0(n1842), .B1(n1798), .Y(n1840) );
  NAND3X1 U3084 ( .A(n1843), .B(n1844), .C(\MEM_CTL/BUS629[1] ), .Y(n1798) );
  CLKINVX1 U3085 ( .A(din[8]), .Y(n1842) );
  NAND3X1 U3086 ( .A(n1844), .B(n1845), .C(n1843), .Y(n1796) );
  CLKINVX1 U3087 ( .A(n1793), .Y(n1843) );
  CLKINVX1 U3088 ( .A(din[24]), .Y(n1841) );
  OAI31X1 U3089 ( .A0(n1844), .A1(\MEM_CTL/BUS629[1] ), .A2(n1793), .B0(n1838), 
        .Y(n1789) );
  NAND2X1 U3090 ( .A(n1827), .B(n1845), .Y(n1838) );
  OAI31X1 U3091 ( .A0(n1844), .A1(n1793), .A2(n1845), .B0(n1837), .Y(n1792) );
  AOI21X1 U3092 ( .A0(\MEM_CTL/BUS629[1] ), .A1(n1827), .B0(n1828), .Y(n1837)
         );
  NOR3X1 U3093 ( .A(n277), .B(n278), .C(n43), .Y(n1828) );
  NOR2X1 U3094 ( .A(n2), .B(n279), .Y(n1827) );
  CLKINVX1 U3095 ( .A(\MEM_CTL/BUS629[1] ), .Y(n1845) );
  AOI31X1 U3096 ( .A0(n277), .A1(n2), .A2(n279), .B0(n1835), .Y(n1793) );
  NOR3X1 U3097 ( .A(n2), .B(n277), .C(n43), .Y(n1835) );
  CLKINVX1 U3098 ( .A(\MEM_CTL/BUS629[0] ), .Y(n1844) );
  CLKINVX1 U3099 ( .A(n1586), .Y(BUS15471[9]) );
  MXI2X1 U3100 ( .A(BUS422[9]), .B(n1846), .S0(NET457), .Y(n1586) );
  OR2X1 U3101 ( .A(BUS7772[9]), .B(cop_dout[9]), .Y(n1846) );
  CLKINVX1 U3102 ( .A(n1588), .Y(BUS15471[8]) );
  MXI2X1 U3103 ( .A(BUS422[8]), .B(n1847), .S0(NET457), .Y(n1588) );
  OR2X1 U3104 ( .A(BUS7772[8]), .B(cop_dout[8]), .Y(n1847) );
  CLKINVX1 U3105 ( .A(n719), .Y(BUS15471[7]) );
  MXI2X1 U3106 ( .A(BUS422[7]), .B(n1848), .S0(NET457), .Y(n719) );
  OR2X1 U3107 ( .A(BUS7772[7]), .B(cop_dout[7]), .Y(n1848) );
  CLKINVX1 U3108 ( .A(n722), .Y(BUS15471[6]) );
  MXI2X1 U3109 ( .A(BUS422[6]), .B(n1849), .S0(NET457), .Y(n722) );
  OR2X1 U3110 ( .A(BUS7772[6]), .B(cop_dout[6]), .Y(n1849) );
  CLKINVX1 U3111 ( .A(n725), .Y(BUS15471[5]) );
  MXI2X1 U3112 ( .A(BUS422[5]), .B(n1850), .S0(NET457), .Y(n725) );
  OR2X1 U3113 ( .A(BUS7772[5]), .B(cop_dout[5]), .Y(n1850) );
  CLKINVX1 U3114 ( .A(n728), .Y(BUS15471[4]) );
  MXI2X1 U3115 ( .A(BUS422[4]), .B(n1851), .S0(NET457), .Y(n728) );
  OR2X1 U3116 ( .A(BUS7772[4]), .B(cop_dout[4]), .Y(n1851) );
  CLKINVX1 U3117 ( .A(n731), .Y(BUS15471[3]) );
  MXI2X1 U3118 ( .A(BUS422[3]), .B(n1852), .S0(NET457), .Y(n731) );
  OR2X1 U3119 ( .A(BUS7772[3]), .B(cop_dout[3]), .Y(n1852) );
  CLKINVX1 U3120 ( .A(n1590), .Y(BUS15471[31]) );
  MXI2X1 U3121 ( .A(BUS422[31]), .B(n1853), .S0(NET457), .Y(n1590) );
  OR2X1 U3122 ( .A(BUS7772[31]), .B(cop_dout[31]), .Y(n1853) );
  CLKINVX1 U3123 ( .A(n1592), .Y(BUS15471[30]) );
  MXI2X1 U3124 ( .A(BUS422[30]), .B(n1854), .S0(NET457), .Y(n1592) );
  OR2X1 U3125 ( .A(BUS7772[30]), .B(cop_dout[30]), .Y(n1854) );
  CLKINVX1 U3126 ( .A(n734), .Y(BUS15471[2]) );
  MXI2X1 U3127 ( .A(BUS422[2]), .B(n1855), .S0(NET457), .Y(n734) );
  OR2X1 U3128 ( .A(BUS7772[2]), .B(cop_dout[2]), .Y(n1855) );
  CLKINVX1 U3129 ( .A(n1594), .Y(BUS15471[29]) );
  MXI2X1 U3130 ( .A(BUS422[29]), .B(n1856), .S0(NET457), .Y(n1594) );
  OR2X1 U3131 ( .A(BUS7772[29]), .B(cop_dout[29]), .Y(n1856) );
  CLKINVX1 U3132 ( .A(n1596), .Y(BUS15471[28]) );
  MXI2X1 U3133 ( .A(BUS422[28]), .B(n1857), .S0(NET457), .Y(n1596) );
  OR2X1 U3134 ( .A(BUS7772[28]), .B(cop_dout[28]), .Y(n1857) );
  CLKINVX1 U3135 ( .A(n1598), .Y(BUS15471[27]) );
  MXI2X1 U3136 ( .A(BUS422[27]), .B(n1858), .S0(NET457), .Y(n1598) );
  OR2X1 U3137 ( .A(BUS7772[27]), .B(cop_dout[27]), .Y(n1858) );
  CLKINVX1 U3138 ( .A(n1600), .Y(BUS15471[26]) );
  MXI2X1 U3139 ( .A(BUS422[26]), .B(n1859), .S0(NET457), .Y(n1600) );
  OR2X1 U3140 ( .A(BUS7772[26]), .B(cop_dout[26]), .Y(n1859) );
  CLKINVX1 U3141 ( .A(n1602), .Y(BUS15471[25]) );
  MXI2X1 U3142 ( .A(BUS422[25]), .B(n1860), .S0(NET457), .Y(n1602) );
  OR2X1 U3143 ( .A(BUS7772[25]), .B(cop_dout[25]), .Y(n1860) );
  CLKINVX1 U3144 ( .A(n1604), .Y(BUS15471[24]) );
  MXI2X1 U3145 ( .A(BUS422[24]), .B(n1861), .S0(NET457), .Y(n1604) );
  OR2X1 U3146 ( .A(BUS7772[24]), .B(cop_dout[24]), .Y(n1861) );
  CLKINVX1 U3147 ( .A(n1606), .Y(BUS15471[23]) );
  MXI2X1 U3148 ( .A(BUS422[23]), .B(n1862), .S0(NET457), .Y(n1606) );
  OR2X1 U3149 ( .A(BUS7772[23]), .B(cop_dout[23]), .Y(n1862) );
  CLKINVX1 U3150 ( .A(n1608), .Y(BUS15471[22]) );
  MXI2X1 U3151 ( .A(BUS422[22]), .B(n1863), .S0(NET457), .Y(n1608) );
  OR2X1 U3152 ( .A(BUS7772[22]), .B(cop_dout[22]), .Y(n1863) );
  CLKINVX1 U3153 ( .A(n1610), .Y(BUS15471[21]) );
  MXI2X1 U3154 ( .A(BUS422[21]), .B(n1864), .S0(NET457), .Y(n1610) );
  OR2X1 U3155 ( .A(BUS7772[21]), .B(cop_dout[21]), .Y(n1864) );
  CLKINVX1 U3156 ( .A(n1612), .Y(BUS15471[20]) );
  MXI2X1 U3157 ( .A(BUS422[20]), .B(n1865), .S0(NET457), .Y(n1612) );
  OR2X1 U3158 ( .A(BUS7772[20]), .B(cop_dout[20]), .Y(n1865) );
  CLKINVX1 U3159 ( .A(n713), .Y(BUS15471[1]) );
  MXI2X1 U3160 ( .A(BUS422[1]), .B(n1866), .S0(NET457), .Y(n713) );
  OR2X1 U3161 ( .A(BUS7772[1]), .B(cop_dout[1]), .Y(n1866) );
  CLKINVX1 U3162 ( .A(n1614), .Y(BUS15471[19]) );
  MXI2X1 U3163 ( .A(BUS422[19]), .B(n1867), .S0(NET457), .Y(n1614) );
  OR2X1 U3164 ( .A(BUS7772[19]), .B(cop_dout[19]), .Y(n1867) );
  CLKINVX1 U3165 ( .A(n1616), .Y(BUS15471[18]) );
  MXI2X1 U3166 ( .A(BUS422[18]), .B(n1868), .S0(NET457), .Y(n1616) );
  OR2X1 U3167 ( .A(BUS7772[18]), .B(cop_dout[18]), .Y(n1868) );
  CLKINVX1 U3168 ( .A(n1618), .Y(BUS15471[17]) );
  MXI2X1 U3169 ( .A(BUS422[17]), .B(n1869), .S0(NET457), .Y(n1618) );
  OR2X1 U3170 ( .A(BUS7772[17]), .B(cop_dout[17]), .Y(n1869) );
  CLKINVX1 U3171 ( .A(n1620), .Y(BUS15471[16]) );
  MXI2X1 U3172 ( .A(BUS422[16]), .B(n1870), .S0(NET457), .Y(n1620) );
  OR2X1 U3173 ( .A(BUS7772[16]), .B(cop_dout[16]), .Y(n1870) );
  CLKINVX1 U3174 ( .A(n1622), .Y(BUS15471[15]) );
  MXI2X1 U3175 ( .A(BUS422[15]), .B(n1871), .S0(NET457), .Y(n1622) );
  OR2X1 U3176 ( .A(BUS7772[15]), .B(cop_dout[15]), .Y(n1871) );
  CLKINVX1 U3177 ( .A(n1624), .Y(BUS15471[14]) );
  MXI2X1 U3178 ( .A(BUS422[14]), .B(n1872), .S0(NET457), .Y(n1624) );
  OR2X1 U3179 ( .A(BUS7772[14]), .B(cop_dout[14]), .Y(n1872) );
  CLKINVX1 U3180 ( .A(n1626), .Y(BUS15471[13]) );
  MXI2X1 U3181 ( .A(BUS422[13]), .B(n1873), .S0(NET457), .Y(n1626) );
  OR2X1 U3182 ( .A(BUS7772[13]), .B(cop_dout[13]), .Y(n1873) );
  CLKINVX1 U3183 ( .A(n1628), .Y(BUS15471[12]) );
  MXI2X1 U3184 ( .A(BUS422[12]), .B(n1874), .S0(NET457), .Y(n1628) );
  OR2X1 U3185 ( .A(BUS7772[12]), .B(cop_dout[12]), .Y(n1874) );
  CLKINVX1 U3186 ( .A(n1630), .Y(BUS15471[11]) );
  MXI2X1 U3187 ( .A(BUS422[11]), .B(n1875), .S0(NET457), .Y(n1630) );
  OR2X1 U3188 ( .A(BUS7772[11]), .B(cop_dout[11]), .Y(n1875) );
  CLKINVX1 U3189 ( .A(n1632), .Y(BUS15471[10]) );
  MXI2X1 U3190 ( .A(BUS422[10]), .B(n1876), .S0(NET457), .Y(n1632) );
  OR2X1 U3191 ( .A(BUS7772[10]), .B(cop_dout[10]), .Y(n1876) );
  CLKINVX1 U3192 ( .A(n737), .Y(BUS15471[0]) );
  MXI2X1 U3193 ( .A(BUS422[0]), .B(n1877), .S0(NET457), .Y(n737) );
  OR2X1 U3194 ( .A(BUS7772[0]), .B(cop_dout[0]), .Y(n1877) );
endmodule

